module main(clk, rst, aes_key, aes_plaintext, reset, aes_ciphertext, ready);
    input clk;
    input rst;
    input[127:0] aes_key;
    input[127:0] aes_plaintext;
    input reset;
    output[127:0] aes_ciphertext;
    output ready;

    reg[7:0] mem_0[255:0]; //tmp4
    reg[7:0] mem_2[255:0]; //tmp6
    reg[7:0] mem_3[255:0]; //tmp7
    reg[7:0] mem_4[255:0]; //tmp8
    reg[7:0] mem_9[255:0]; //tmp4
    reg[7:0] mem_10[255:0]; //tmp4
    reg[7:0] mem_11[255:0]; //tmp4
    reg[7:0] mem_12[255:0]; //tmp4
    reg[7:0] mem_13[255:0]; //tmp4
    reg[7:0] mem_14[255:0]; //tmp4
    reg[7:0] mem_15[255:0]; //tmp4
    reg[7:0] mem_16[255:0]; //tmp4
    reg[7:0] mem_17[255:0]; //tmp4
    reg[7:0] mem_18[255:0]; //tmp4
    reg[7:0] mem_19[255:0]; //tmp4
    reg[7:0] mem_20[255:0]; //tmp4
    reg[7:0] mem_21[255:0]; //tmp4
    reg[7:0] mem_22[255:0]; //tmp4
    reg[7:0] mem_23[255:0]; //tmp4
    reg[7:0] mem_24[255:0]; //tmp7
    reg[7:0] mem_25[255:0]; //tmp8
    reg[7:0] mem_26[255:0]; //tmp7
    reg[7:0] mem_27[255:0]; //tmp8
    reg[7:0] mem_28[255:0]; //tmp7
    reg[7:0] mem_29[255:0]; //tmp8
    reg[7:0] mem_30[255:0]; //tmp7
    reg[7:0] mem_31[255:0]; //tmp8
    reg[7:0] mem_32[255:0]; //tmp7
    reg[7:0] mem_33[255:0]; //tmp8
    reg[7:0] mem_34[255:0]; //tmp7
    reg[7:0] mem_35[255:0]; //tmp8
    reg[7:0] mem_36[255:0]; //tmp7
    reg[7:0] mem_37[255:0]; //tmp8
    reg[7:0] mem_38[255:0]; //tmp7
    reg[7:0] mem_39[255:0]; //tmp8
    reg[7:0] mem_40[255:0]; //tmp7
    reg[7:0] mem_41[255:0]; //tmp8
    reg[7:0] mem_42[255:0]; //tmp7
    reg[7:0] mem_43[255:0]; //tmp8
    reg[7:0] mem_44[255:0]; //tmp7
    reg[7:0] mem_45[255:0]; //tmp8
    reg[7:0] mem_46[255:0]; //tmp7
    reg[7:0] mem_47[255:0]; //tmp8
    reg[7:0] mem_48[255:0]; //tmp7
    reg[7:0] mem_49[255:0]; //tmp8
    reg[7:0] mem_50[255:0]; //tmp7
    reg[7:0] mem_51[255:0]; //tmp8
    reg[7:0] mem_52[255:0]; //tmp7
    reg[7:0] mem_53[255:0]; //tmp8
    reg[7:0] mem_54[255:0]; //tmp4
    reg[7:0] mem_55[255:0]; //tmp4
    reg[7:0] mem_56[255:0]; //tmp4
    reg[7:0] mem_57[255:0]; //tmp4
    reg[3:0] counter;
    reg[127:0] tmp0;
    reg[127:0] tmp1;

    wire const_0_1;
    wire const_1_0;
    wire const_2_0;
    wire const_3_1;
    wire[3:0] const_4_0;
    wire[3:0] const_5_10;
    wire const_6_1;
    wire const_7_0;
    wire[3:0] const_8_9;
    wire const_9_0;
    wire const_10_0;
    wire const_11_0;
    wire const_12_0;
    wire const_13_0;
    wire const_14_0;
    wire[3:0] const_15_10;
    wire[7:0] tmp13;
    wire[7:0] tmp14;
    wire[7:0] tmp15;
    wire[7:0] tmp16;
    wire[7:0] tmp17;
    wire[7:0] tmp18;
    wire[7:0] tmp19;
    wire[7:0] tmp20;
    wire[7:0] tmp21;
    wire[7:0] tmp22;
    wire[7:0] tmp23;
    wire[7:0] tmp24;
    wire[7:0] tmp25;
    wire[7:0] tmp26;
    wire[7:0] tmp27;
    wire[7:0] tmp28;
    wire[7:0] tmp29;
    wire[7:0] tmp30;
    wire[7:0] tmp31;
    wire[7:0] tmp32;
    wire[7:0] tmp33;
    wire[7:0] tmp34;
    wire[7:0] tmp35;
    wire[7:0] tmp36;
    wire[7:0] tmp37;
    wire[7:0] tmp38;
    wire[7:0] tmp39;
    wire[7:0] tmp40;
    wire[7:0] tmp41;
    wire[7:0] tmp42;
    wire[7:0] tmp43;
    wire[7:0] tmp44;
    wire[127:0] tmp45;
    wire[7:0] tmp46;
    wire[7:0] tmp47;
    wire[7:0] tmp48;
    wire[7:0] tmp49;
    wire[7:0] tmp50;
    wire[7:0] tmp51;
    wire[7:0] tmp52;
    wire[7:0] tmp53;
    wire[7:0] tmp54;
    wire[7:0] tmp55;
    wire[7:0] tmp56;
    wire[7:0] tmp57;
    wire[7:0] tmp58;
    wire[7:0] tmp59;
    wire[7:0] tmp60;
    wire[7:0] tmp61;
    wire[127:0] tmp62;
    wire[31:0] tmp63;
    wire[31:0] tmp64;
    wire[31:0] tmp65;
    wire[31:0] tmp66;
    wire[7:0] tmp67;
    wire[7:0] tmp68;
    wire[7:0] tmp69;
    wire[7:0] tmp70;
    wire[7:0] tmp71;
    wire[7:0] tmp72;
    wire[7:0] tmp73;
    wire[7:0] tmp74;
    wire[7:0] tmp75;
    wire[7:0] tmp76;
    wire[7:0] tmp77;
    wire[7:0] tmp78;
    wire[7:0] tmp79;
    wire[7:0] tmp80;
    wire[7:0] tmp81;
    wire[7:0] tmp82;
    wire[7:0] tmp83;
    wire[7:0] tmp84;
    wire[7:0] tmp85;
    wire[7:0] tmp86;
    wire[7:0] tmp87;
    wire[7:0] tmp88;
    wire[7:0] tmp89;
    wire[7:0] tmp90;
    wire[31:0] tmp91;
    wire[7:0] tmp92;
    wire[7:0] tmp93;
    wire[7:0] tmp94;
    wire[7:0] tmp95;
    wire[7:0] tmp96;
    wire[7:0] tmp97;
    wire[7:0] tmp98;
    wire[7:0] tmp99;
    wire[7:0] tmp100;
    wire[7:0] tmp101;
    wire[7:0] tmp102;
    wire[7:0] tmp103;
    wire[7:0] tmp104;
    wire[7:0] tmp105;
    wire[7:0] tmp106;
    wire[7:0] tmp107;
    wire[7:0] tmp108;
    wire[7:0] tmp109;
    wire[7:0] tmp110;
    wire[7:0] tmp111;
    wire[7:0] tmp112;
    wire[7:0] tmp113;
    wire[7:0] tmp114;
    wire[7:0] tmp115;
    wire[31:0] tmp116;
    wire[7:0] tmp117;
    wire[7:0] tmp118;
    wire[7:0] tmp119;
    wire[7:0] tmp120;
    wire[7:0] tmp121;
    wire[7:0] tmp122;
    wire[7:0] tmp123;
    wire[7:0] tmp124;
    wire[7:0] tmp125;
    wire[7:0] tmp126;
    wire[7:0] tmp127;
    wire[7:0] tmp128;
    wire[7:0] tmp129;
    wire[7:0] tmp130;
    wire[7:0] tmp131;
    wire[7:0] tmp132;
    wire[7:0] tmp133;
    wire[7:0] tmp134;
    wire[7:0] tmp135;
    wire[7:0] tmp136;
    wire[7:0] tmp137;
    wire[7:0] tmp138;
    wire[7:0] tmp139;
    wire[7:0] tmp140;
    wire[31:0] tmp141;
    wire[7:0] tmp142;
    wire[7:0] tmp143;
    wire[7:0] tmp144;
    wire[7:0] tmp145;
    wire[7:0] tmp146;
    wire[7:0] tmp147;
    wire[7:0] tmp148;
    wire[7:0] tmp149;
    wire[7:0] tmp150;
    wire[7:0] tmp151;
    wire[7:0] tmp152;
    wire[7:0] tmp153;
    wire[7:0] tmp154;
    wire[7:0] tmp155;
    wire[7:0] tmp156;
    wire[7:0] tmp157;
    wire[7:0] tmp158;
    wire[7:0] tmp159;
    wire[7:0] tmp160;
    wire[7:0] tmp161;
    wire[7:0] tmp162;
    wire[7:0] tmp163;
    wire[7:0] tmp164;
    wire[7:0] tmp165;
    wire[31:0] tmp166;
    wire[127:0] tmp167;
    wire[31:0] tmp168;
    wire[31:0] tmp169;
    wire[31:0] tmp170;
    wire[31:0] tmp171;
    wire[7:0] tmp172;
    wire[7:0] tmp173;
    wire[7:0] tmp174;
    wire[7:0] tmp175;
    wire[3:0] tmp179;
    wire[7:0] tmp180;
    wire[7:0] tmp181;
    wire[7:0] tmp182;
    wire[7:0] tmp183;
    wire[7:0] tmp184;
    wire[7:0] tmp185;
    wire[7:0] tmp186;
    wire[31:0] tmp187;
    wire[31:0] tmp188;
    wire[31:0] tmp189;
    wire[31:0] tmp190;
    wire[31:0] tmp191;
    wire[127:0] tmp192;
    wire[127:0] tmp193;
    wire tmp194;
    wire tmp195;
    wire tmp197;
    wire[2:0] tmp200;
    wire[3:0] tmp201;
    wire[3:0] tmp202;
    wire tmp212;
    wire tmp215;
    wire tmp218;
    wire tmp219;
    wire tmp221;
    wire tmp223;
    wire tmp224;
    wire[3:0] tmp226;
    wire[3:0] tmp227;
    wire[3:0] tmp228;
    wire[3:0] tmp229;
    wire[126:0] tmp230;
    wire[127:0] tmp232;
    wire[127:0] tmp233;
    wire[127:0] tmp234;
    wire[127:0] tmp235;
    wire[127:0] tmp236;
    wire[127:0] tmp237;
    wire[127:0] tmp238;
    wire[127:0] tmp240;
    wire[127:0] tmp241;
    wire[127:0] tmp242;
    wire[127:0] tmp243;

    initial begin
        mem_0[0]=8'h63;
        mem_0[1]=8'h7c;
        mem_0[2]=8'h77;
        mem_0[3]=8'h7b;
        mem_0[4]=8'hf2;
        mem_0[5]=8'h6b;
        mem_0[6]=8'h6f;
        mem_0[7]=8'hc5;
        mem_0[8]=8'h30;
        mem_0[9]=8'h1;
        mem_0[10]=8'h67;
        mem_0[11]=8'h2b;
        mem_0[12]=8'hfe;
        mem_0[13]=8'hd7;
        mem_0[14]=8'hab;
        mem_0[15]=8'h76;
        mem_0[16]=8'hca;
        mem_0[17]=8'h82;
        mem_0[18]=8'hc9;
        mem_0[19]=8'h7d;
        mem_0[20]=8'hfa;
        mem_0[21]=8'h59;
        mem_0[22]=8'h47;
        mem_0[23]=8'hf0;
        mem_0[24]=8'had;
        mem_0[25]=8'hd4;
        mem_0[26]=8'ha2;
        mem_0[27]=8'haf;
        mem_0[28]=8'h9c;
        mem_0[29]=8'ha4;
        mem_0[30]=8'h72;
        mem_0[31]=8'hc0;
        mem_0[32]=8'hb7;
        mem_0[33]=8'hfd;
        mem_0[34]=8'h93;
        mem_0[35]=8'h26;
        mem_0[36]=8'h36;
        mem_0[37]=8'h3f;
        mem_0[38]=8'hf7;
        mem_0[39]=8'hcc;
        mem_0[40]=8'h34;
        mem_0[41]=8'ha5;
        mem_0[42]=8'he5;
        mem_0[43]=8'hf1;
        mem_0[44]=8'h71;
        mem_0[45]=8'hd8;
        mem_0[46]=8'h31;
        mem_0[47]=8'h15;
        mem_0[48]=8'h4;
        mem_0[49]=8'hc7;
        mem_0[50]=8'h23;
        mem_0[51]=8'hc3;
        mem_0[52]=8'h18;
        mem_0[53]=8'h96;
        mem_0[54]=8'h5;
        mem_0[55]=8'h9a;
        mem_0[56]=8'h7;
        mem_0[57]=8'h12;
        mem_0[58]=8'h80;
        mem_0[59]=8'he2;
        mem_0[60]=8'heb;
        mem_0[61]=8'h27;
        mem_0[62]=8'hb2;
        mem_0[63]=8'h75;
        mem_0[64]=8'h9;
        mem_0[65]=8'h83;
        mem_0[66]=8'h2c;
        mem_0[67]=8'h1a;
        mem_0[68]=8'h1b;
        mem_0[69]=8'h6e;
        mem_0[70]=8'h5a;
        mem_0[71]=8'ha0;
        mem_0[72]=8'h52;
        mem_0[73]=8'h3b;
        mem_0[74]=8'hd6;
        mem_0[75]=8'hb3;
        mem_0[76]=8'h29;
        mem_0[77]=8'he3;
        mem_0[78]=8'h2f;
        mem_0[79]=8'h84;
        mem_0[80]=8'h53;
        mem_0[81]=8'hd1;
        mem_0[82]=8'h0;
        mem_0[83]=8'hed;
        mem_0[84]=8'h20;
        mem_0[85]=8'hfc;
        mem_0[86]=8'hb1;
        mem_0[87]=8'h5b;
        mem_0[88]=8'h6a;
        mem_0[89]=8'hcb;
        mem_0[90]=8'hbe;
        mem_0[91]=8'h39;
        mem_0[92]=8'h4a;
        mem_0[93]=8'h4c;
        mem_0[94]=8'h58;
        mem_0[95]=8'hcf;
        mem_0[96]=8'hd0;
        mem_0[97]=8'hef;
        mem_0[98]=8'haa;
        mem_0[99]=8'hfb;
        mem_0[100]=8'h43;
        mem_0[101]=8'h4d;
        mem_0[102]=8'h33;
        mem_0[103]=8'h85;
        mem_0[104]=8'h45;
        mem_0[105]=8'hf9;
        mem_0[106]=8'h2;
        mem_0[107]=8'h7f;
        mem_0[108]=8'h50;
        mem_0[109]=8'h3c;
        mem_0[110]=8'h9f;
        mem_0[111]=8'ha8;
        mem_0[112]=8'h51;
        mem_0[113]=8'ha3;
        mem_0[114]=8'h40;
        mem_0[115]=8'h8f;
        mem_0[116]=8'h92;
        mem_0[117]=8'h9d;
        mem_0[118]=8'h38;
        mem_0[119]=8'hf5;
        mem_0[120]=8'hbc;
        mem_0[121]=8'hb6;
        mem_0[122]=8'hda;
        mem_0[123]=8'h21;
        mem_0[124]=8'h10;
        mem_0[125]=8'hff;
        mem_0[126]=8'hf3;
        mem_0[127]=8'hd2;
        mem_0[128]=8'hcd;
        mem_0[129]=8'hc;
        mem_0[130]=8'h13;
        mem_0[131]=8'hec;
        mem_0[132]=8'h5f;
        mem_0[133]=8'h97;
        mem_0[134]=8'h44;
        mem_0[135]=8'h17;
        mem_0[136]=8'hc4;
        mem_0[137]=8'ha7;
        mem_0[138]=8'h7e;
        mem_0[139]=8'h3d;
        mem_0[140]=8'h64;
        mem_0[141]=8'h5d;
        mem_0[142]=8'h19;
        mem_0[143]=8'h73;
        mem_0[144]=8'h60;
        mem_0[145]=8'h81;
        mem_0[146]=8'h4f;
        mem_0[147]=8'hdc;
        mem_0[148]=8'h22;
        mem_0[149]=8'h2a;
        mem_0[150]=8'h90;
        mem_0[151]=8'h88;
        mem_0[152]=8'h46;
        mem_0[153]=8'hee;
        mem_0[154]=8'hb8;
        mem_0[155]=8'h14;
        mem_0[156]=8'hde;
        mem_0[157]=8'h5e;
        mem_0[158]=8'hb;
        mem_0[159]=8'hdb;
        mem_0[160]=8'he0;
        mem_0[161]=8'h32;
        mem_0[162]=8'h3a;
        mem_0[163]=8'ha;
        mem_0[164]=8'h49;
        mem_0[165]=8'h6;
        mem_0[166]=8'h24;
        mem_0[167]=8'h5c;
        mem_0[168]=8'hc2;
        mem_0[169]=8'hd3;
        mem_0[170]=8'hac;
        mem_0[171]=8'h62;
        mem_0[172]=8'h91;
        mem_0[173]=8'h95;
        mem_0[174]=8'he4;
        mem_0[175]=8'h79;
        mem_0[176]=8'he7;
        mem_0[177]=8'hc8;
        mem_0[178]=8'h37;
        mem_0[179]=8'h6d;
        mem_0[180]=8'h8d;
        mem_0[181]=8'hd5;
        mem_0[182]=8'h4e;
        mem_0[183]=8'ha9;
        mem_0[184]=8'h6c;
        mem_0[185]=8'h56;
        mem_0[186]=8'hf4;
        mem_0[187]=8'hea;
        mem_0[188]=8'h65;
        mem_0[189]=8'h7a;
        mem_0[190]=8'hae;
        mem_0[191]=8'h8;
        mem_0[192]=8'hba;
        mem_0[193]=8'h78;
        mem_0[194]=8'h25;
        mem_0[195]=8'h2e;
        mem_0[196]=8'h1c;
        mem_0[197]=8'ha6;
        mem_0[198]=8'hb4;
        mem_0[199]=8'hc6;
        mem_0[200]=8'he8;
        mem_0[201]=8'hdd;
        mem_0[202]=8'h74;
        mem_0[203]=8'h1f;
        mem_0[204]=8'h4b;
        mem_0[205]=8'hbd;
        mem_0[206]=8'h8b;
        mem_0[207]=8'h8a;
        mem_0[208]=8'h70;
        mem_0[209]=8'h3e;
        mem_0[210]=8'hb5;
        mem_0[211]=8'h66;
        mem_0[212]=8'h48;
        mem_0[213]=8'h3;
        mem_0[214]=8'hf6;
        mem_0[215]=8'he;
        mem_0[216]=8'h61;
        mem_0[217]=8'h35;
        mem_0[218]=8'h57;
        mem_0[219]=8'hb9;
        mem_0[220]=8'h86;
        mem_0[221]=8'hc1;
        mem_0[222]=8'h1d;
        mem_0[223]=8'h9e;
        mem_0[224]=8'he1;
        mem_0[225]=8'hf8;
        mem_0[226]=8'h98;
        mem_0[227]=8'h11;
        mem_0[228]=8'h69;
        mem_0[229]=8'hd9;
        mem_0[230]=8'h8e;
        mem_0[231]=8'h94;
        mem_0[232]=8'h9b;
        mem_0[233]=8'h1e;
        mem_0[234]=8'h87;
        mem_0[235]=8'he9;
        mem_0[236]=8'hce;
        mem_0[237]=8'h55;
        mem_0[238]=8'h28;
        mem_0[239]=8'hdf;
        mem_0[240]=8'h8c;
        mem_0[241]=8'ha1;
        mem_0[242]=8'h89;
        mem_0[243]=8'hd;
        mem_0[244]=8'hbf;
        mem_0[245]=8'he6;
        mem_0[246]=8'h42;
        mem_0[247]=8'h68;
        mem_0[248]=8'h41;
        mem_0[249]=8'h99;
        mem_0[250]=8'h2d;
        mem_0[251]=8'hf;
        mem_0[252]=8'hb0;
        mem_0[253]=8'h54;
        mem_0[254]=8'hbb;
        mem_0[255]=8'h16;
    end

    initial begin
        mem_2[0]=8'h8d;
        mem_2[1]=8'h1;
        mem_2[2]=8'h2;
        mem_2[3]=8'h4;
        mem_2[4]=8'h8;
        mem_2[5]=8'h10;
        mem_2[6]=8'h20;
        mem_2[7]=8'h40;
        mem_2[8]=8'h80;
        mem_2[9]=8'h1b;
        mem_2[10]=8'h36;
        mem_2[11]=8'h6c;
        mem_2[12]=8'hd8;
        mem_2[13]=8'hab;
        mem_2[14]=8'h4d;
        mem_2[15]=8'h9a;
        mem_2[16]=8'h2f;
        mem_2[17]=8'h5e;
        mem_2[18]=8'hbc;
        mem_2[19]=8'h63;
        mem_2[20]=8'hc6;
        mem_2[21]=8'h97;
        mem_2[22]=8'h35;
        mem_2[23]=8'h6a;
        mem_2[24]=8'hd4;
        mem_2[25]=8'hb3;
        mem_2[26]=8'h7d;
        mem_2[27]=8'hfa;
        mem_2[28]=8'hef;
        mem_2[29]=8'hc5;
        mem_2[30]=8'h91;
        mem_2[31]=8'h39;
        mem_2[32]=8'h72;
        mem_2[33]=8'he4;
        mem_2[34]=8'hd3;
        mem_2[35]=8'hbd;
        mem_2[36]=8'h61;
        mem_2[37]=8'hc2;
        mem_2[38]=8'h9f;
        mem_2[39]=8'h25;
        mem_2[40]=8'h4a;
        mem_2[41]=8'h94;
        mem_2[42]=8'h33;
        mem_2[43]=8'h66;
        mem_2[44]=8'hcc;
        mem_2[45]=8'h83;
        mem_2[46]=8'h1d;
        mem_2[47]=8'h3a;
        mem_2[48]=8'h74;
        mem_2[49]=8'he8;
        mem_2[50]=8'hcb;
        mem_2[51]=8'h8d;
        mem_2[52]=8'h1;
        mem_2[53]=8'h2;
        mem_2[54]=8'h4;
        mem_2[55]=8'h8;
        mem_2[56]=8'h10;
        mem_2[57]=8'h20;
        mem_2[58]=8'h40;
        mem_2[59]=8'h80;
        mem_2[60]=8'h1b;
        mem_2[61]=8'h36;
        mem_2[62]=8'h6c;
        mem_2[63]=8'hd8;
        mem_2[64]=8'hab;
        mem_2[65]=8'h4d;
        mem_2[66]=8'h9a;
        mem_2[67]=8'h2f;
        mem_2[68]=8'h5e;
        mem_2[69]=8'hbc;
        mem_2[70]=8'h63;
        mem_2[71]=8'hc6;
        mem_2[72]=8'h97;
        mem_2[73]=8'h35;
        mem_2[74]=8'h6a;
        mem_2[75]=8'hd4;
        mem_2[76]=8'hb3;
        mem_2[77]=8'h7d;
        mem_2[78]=8'hfa;
        mem_2[79]=8'hef;
        mem_2[80]=8'hc5;
        mem_2[81]=8'h91;
        mem_2[82]=8'h39;
        mem_2[83]=8'h72;
        mem_2[84]=8'he4;
        mem_2[85]=8'hd3;
        mem_2[86]=8'hbd;
        mem_2[87]=8'h61;
        mem_2[88]=8'hc2;
        mem_2[89]=8'h9f;
        mem_2[90]=8'h25;
        mem_2[91]=8'h4a;
        mem_2[92]=8'h94;
        mem_2[93]=8'h33;
        mem_2[94]=8'h66;
        mem_2[95]=8'hcc;
        mem_2[96]=8'h83;
        mem_2[97]=8'h1d;
        mem_2[98]=8'h3a;
        mem_2[99]=8'h74;
        mem_2[100]=8'he8;
        mem_2[101]=8'hcb;
        mem_2[102]=8'h8d;
        mem_2[103]=8'h1;
        mem_2[104]=8'h2;
        mem_2[105]=8'h4;
        mem_2[106]=8'h8;
        mem_2[107]=8'h10;
        mem_2[108]=8'h20;
        mem_2[109]=8'h40;
        mem_2[110]=8'h80;
        mem_2[111]=8'h1b;
        mem_2[112]=8'h36;
        mem_2[113]=8'h6c;
        mem_2[114]=8'hd8;
        mem_2[115]=8'hab;
        mem_2[116]=8'h4d;
        mem_2[117]=8'h9a;
        mem_2[118]=8'h2f;
        mem_2[119]=8'h5e;
        mem_2[120]=8'hbc;
        mem_2[121]=8'h63;
        mem_2[122]=8'hc6;
        mem_2[123]=8'h97;
        mem_2[124]=8'h35;
        mem_2[125]=8'h6a;
        mem_2[126]=8'hd4;
        mem_2[127]=8'hb3;
        mem_2[128]=8'h7d;
        mem_2[129]=8'hfa;
        mem_2[130]=8'hef;
        mem_2[131]=8'hc5;
        mem_2[132]=8'h91;
        mem_2[133]=8'h39;
        mem_2[134]=8'h72;
        mem_2[135]=8'he4;
        mem_2[136]=8'hd3;
        mem_2[137]=8'hbd;
        mem_2[138]=8'h61;
        mem_2[139]=8'hc2;
        mem_2[140]=8'h9f;
        mem_2[141]=8'h25;
        mem_2[142]=8'h4a;
        mem_2[143]=8'h94;
        mem_2[144]=8'h33;
        mem_2[145]=8'h66;
        mem_2[146]=8'hcc;
        mem_2[147]=8'h83;
        mem_2[148]=8'h1d;
        mem_2[149]=8'h3a;
        mem_2[150]=8'h74;
        mem_2[151]=8'he8;
        mem_2[152]=8'hcb;
        mem_2[153]=8'h8d;
        mem_2[154]=8'h1;
        mem_2[155]=8'h2;
        mem_2[156]=8'h4;
        mem_2[157]=8'h8;
        mem_2[158]=8'h10;
        mem_2[159]=8'h20;
        mem_2[160]=8'h40;
        mem_2[161]=8'h80;
        mem_2[162]=8'h1b;
        mem_2[163]=8'h36;
        mem_2[164]=8'h6c;
        mem_2[165]=8'hd8;
        mem_2[166]=8'hab;
        mem_2[167]=8'h4d;
        mem_2[168]=8'h9a;
        mem_2[169]=8'h2f;
        mem_2[170]=8'h5e;
        mem_2[171]=8'hbc;
        mem_2[172]=8'h63;
        mem_2[173]=8'hc6;
        mem_2[174]=8'h97;
        mem_2[175]=8'h35;
        mem_2[176]=8'h6a;
        mem_2[177]=8'hd4;
        mem_2[178]=8'hb3;
        mem_2[179]=8'h7d;
        mem_2[180]=8'hfa;
        mem_2[181]=8'hef;
        mem_2[182]=8'hc5;
        mem_2[183]=8'h91;
        mem_2[184]=8'h39;
        mem_2[185]=8'h72;
        mem_2[186]=8'he4;
        mem_2[187]=8'hd3;
        mem_2[188]=8'hbd;
        mem_2[189]=8'h61;
        mem_2[190]=8'hc2;
        mem_2[191]=8'h9f;
        mem_2[192]=8'h25;
        mem_2[193]=8'h4a;
        mem_2[194]=8'h94;
        mem_2[195]=8'h33;
        mem_2[196]=8'h66;
        mem_2[197]=8'hcc;
        mem_2[198]=8'h83;
        mem_2[199]=8'h1d;
        mem_2[200]=8'h3a;
        mem_2[201]=8'h74;
        mem_2[202]=8'he8;
        mem_2[203]=8'hcb;
        mem_2[204]=8'h8d;
        mem_2[205]=8'h1;
        mem_2[206]=8'h2;
        mem_2[207]=8'h4;
        mem_2[208]=8'h8;
        mem_2[209]=8'h10;
        mem_2[210]=8'h20;
        mem_2[211]=8'h40;
        mem_2[212]=8'h80;
        mem_2[213]=8'h1b;
        mem_2[214]=8'h36;
        mem_2[215]=8'h6c;
        mem_2[216]=8'hd8;
        mem_2[217]=8'hab;
        mem_2[218]=8'h4d;
        mem_2[219]=8'h9a;
        mem_2[220]=8'h2f;
        mem_2[221]=8'h5e;
        mem_2[222]=8'hbc;
        mem_2[223]=8'h63;
        mem_2[224]=8'hc6;
        mem_2[225]=8'h97;
        mem_2[226]=8'h35;
        mem_2[227]=8'h6a;
        mem_2[228]=8'hd4;
        mem_2[229]=8'hb3;
        mem_2[230]=8'h7d;
        mem_2[231]=8'hfa;
        mem_2[232]=8'hef;
        mem_2[233]=8'hc5;
        mem_2[234]=8'h91;
        mem_2[235]=8'h39;
        mem_2[236]=8'h72;
        mem_2[237]=8'he4;
        mem_2[238]=8'hd3;
        mem_2[239]=8'hbd;
        mem_2[240]=8'h61;
        mem_2[241]=8'hc2;
        mem_2[242]=8'h9f;
        mem_2[243]=8'h25;
        mem_2[244]=8'h4a;
        mem_2[245]=8'h94;
        mem_2[246]=8'h33;
        mem_2[247]=8'h66;
        mem_2[248]=8'hcc;
        mem_2[249]=8'h83;
        mem_2[250]=8'h1d;
        mem_2[251]=8'h3a;
        mem_2[252]=8'h74;
        mem_2[253]=8'he8;
        mem_2[254]=8'hcb;
        mem_2[255]=8'h8d;
    end

    initial begin
        mem_3[0]=8'h0;
        mem_3[1]=8'h2;
        mem_3[2]=8'h4;
        mem_3[3]=8'h6;
        mem_3[4]=8'h8;
        mem_3[5]=8'ha;
        mem_3[6]=8'hc;
        mem_3[7]=8'he;
        mem_3[8]=8'h10;
        mem_3[9]=8'h12;
        mem_3[10]=8'h14;
        mem_3[11]=8'h16;
        mem_3[12]=8'h18;
        mem_3[13]=8'h1a;
        mem_3[14]=8'h1c;
        mem_3[15]=8'h1e;
        mem_3[16]=8'h20;
        mem_3[17]=8'h22;
        mem_3[18]=8'h24;
        mem_3[19]=8'h26;
        mem_3[20]=8'h28;
        mem_3[21]=8'h2a;
        mem_3[22]=8'h2c;
        mem_3[23]=8'h2e;
        mem_3[24]=8'h30;
        mem_3[25]=8'h32;
        mem_3[26]=8'h34;
        mem_3[27]=8'h36;
        mem_3[28]=8'h38;
        mem_3[29]=8'h3a;
        mem_3[30]=8'h3c;
        mem_3[31]=8'h3e;
        mem_3[32]=8'h40;
        mem_3[33]=8'h42;
        mem_3[34]=8'h44;
        mem_3[35]=8'h46;
        mem_3[36]=8'h48;
        mem_3[37]=8'h4a;
        mem_3[38]=8'h4c;
        mem_3[39]=8'h4e;
        mem_3[40]=8'h50;
        mem_3[41]=8'h52;
        mem_3[42]=8'h54;
        mem_3[43]=8'h56;
        mem_3[44]=8'h58;
        mem_3[45]=8'h5a;
        mem_3[46]=8'h5c;
        mem_3[47]=8'h5e;
        mem_3[48]=8'h60;
        mem_3[49]=8'h62;
        mem_3[50]=8'h64;
        mem_3[51]=8'h66;
        mem_3[52]=8'h68;
        mem_3[53]=8'h6a;
        mem_3[54]=8'h6c;
        mem_3[55]=8'h6e;
        mem_3[56]=8'h70;
        mem_3[57]=8'h72;
        mem_3[58]=8'h74;
        mem_3[59]=8'h76;
        mem_3[60]=8'h78;
        mem_3[61]=8'h7a;
        mem_3[62]=8'h7c;
        mem_3[63]=8'h7e;
        mem_3[64]=8'h80;
        mem_3[65]=8'h82;
        mem_3[66]=8'h84;
        mem_3[67]=8'h86;
        mem_3[68]=8'h88;
        mem_3[69]=8'h8a;
        mem_3[70]=8'h8c;
        mem_3[71]=8'h8e;
        mem_3[72]=8'h90;
        mem_3[73]=8'h92;
        mem_3[74]=8'h94;
        mem_3[75]=8'h96;
        mem_3[76]=8'h98;
        mem_3[77]=8'h9a;
        mem_3[78]=8'h9c;
        mem_3[79]=8'h9e;
        mem_3[80]=8'ha0;
        mem_3[81]=8'ha2;
        mem_3[82]=8'ha4;
        mem_3[83]=8'ha6;
        mem_3[84]=8'ha8;
        mem_3[85]=8'haa;
        mem_3[86]=8'hac;
        mem_3[87]=8'hae;
        mem_3[88]=8'hb0;
        mem_3[89]=8'hb2;
        mem_3[90]=8'hb4;
        mem_3[91]=8'hb6;
        mem_3[92]=8'hb8;
        mem_3[93]=8'hba;
        mem_3[94]=8'hbc;
        mem_3[95]=8'hbe;
        mem_3[96]=8'hc0;
        mem_3[97]=8'hc2;
        mem_3[98]=8'hc4;
        mem_3[99]=8'hc6;
        mem_3[100]=8'hc8;
        mem_3[101]=8'hca;
        mem_3[102]=8'hcc;
        mem_3[103]=8'hce;
        mem_3[104]=8'hd0;
        mem_3[105]=8'hd2;
        mem_3[106]=8'hd4;
        mem_3[107]=8'hd6;
        mem_3[108]=8'hd8;
        mem_3[109]=8'hda;
        mem_3[110]=8'hdc;
        mem_3[111]=8'hde;
        mem_3[112]=8'he0;
        mem_3[113]=8'he2;
        mem_3[114]=8'he4;
        mem_3[115]=8'he6;
        mem_3[116]=8'he8;
        mem_3[117]=8'hea;
        mem_3[118]=8'hec;
        mem_3[119]=8'hee;
        mem_3[120]=8'hf0;
        mem_3[121]=8'hf2;
        mem_3[122]=8'hf4;
        mem_3[123]=8'hf6;
        mem_3[124]=8'hf8;
        mem_3[125]=8'hfa;
        mem_3[126]=8'hfc;
        mem_3[127]=8'hfe;
        mem_3[128]=8'h1b;
        mem_3[129]=8'h19;
        mem_3[130]=8'h1f;
        mem_3[131]=8'h1d;
        mem_3[132]=8'h13;
        mem_3[133]=8'h11;
        mem_3[134]=8'h17;
        mem_3[135]=8'h15;
        mem_3[136]=8'hb;
        mem_3[137]=8'h9;
        mem_3[138]=8'hf;
        mem_3[139]=8'hd;
        mem_3[140]=8'h3;
        mem_3[141]=8'h1;
        mem_3[142]=8'h7;
        mem_3[143]=8'h5;
        mem_3[144]=8'h3b;
        mem_3[145]=8'h39;
        mem_3[146]=8'h3f;
        mem_3[147]=8'h3d;
        mem_3[148]=8'h33;
        mem_3[149]=8'h31;
        mem_3[150]=8'h37;
        mem_3[151]=8'h35;
        mem_3[152]=8'h2b;
        mem_3[153]=8'h29;
        mem_3[154]=8'h2f;
        mem_3[155]=8'h2d;
        mem_3[156]=8'h23;
        mem_3[157]=8'h21;
        mem_3[158]=8'h27;
        mem_3[159]=8'h25;
        mem_3[160]=8'h5b;
        mem_3[161]=8'h59;
        mem_3[162]=8'h5f;
        mem_3[163]=8'h5d;
        mem_3[164]=8'h53;
        mem_3[165]=8'h51;
        mem_3[166]=8'h57;
        mem_3[167]=8'h55;
        mem_3[168]=8'h4b;
        mem_3[169]=8'h49;
        mem_3[170]=8'h4f;
        mem_3[171]=8'h4d;
        mem_3[172]=8'h43;
        mem_3[173]=8'h41;
        mem_3[174]=8'h47;
        mem_3[175]=8'h45;
        mem_3[176]=8'h7b;
        mem_3[177]=8'h79;
        mem_3[178]=8'h7f;
        mem_3[179]=8'h7d;
        mem_3[180]=8'h73;
        mem_3[181]=8'h71;
        mem_3[182]=8'h77;
        mem_3[183]=8'h75;
        mem_3[184]=8'h6b;
        mem_3[185]=8'h69;
        mem_3[186]=8'h6f;
        mem_3[187]=8'h6d;
        mem_3[188]=8'h63;
        mem_3[189]=8'h61;
        mem_3[190]=8'h67;
        mem_3[191]=8'h65;
        mem_3[192]=8'h9b;
        mem_3[193]=8'h99;
        mem_3[194]=8'h9f;
        mem_3[195]=8'h9d;
        mem_3[196]=8'h93;
        mem_3[197]=8'h91;
        mem_3[198]=8'h97;
        mem_3[199]=8'h95;
        mem_3[200]=8'h8b;
        mem_3[201]=8'h89;
        mem_3[202]=8'h8f;
        mem_3[203]=8'h8d;
        mem_3[204]=8'h83;
        mem_3[205]=8'h81;
        mem_3[206]=8'h87;
        mem_3[207]=8'h85;
        mem_3[208]=8'hbb;
        mem_3[209]=8'hb9;
        mem_3[210]=8'hbf;
        mem_3[211]=8'hbd;
        mem_3[212]=8'hb3;
        mem_3[213]=8'hb1;
        mem_3[214]=8'hb7;
        mem_3[215]=8'hb5;
        mem_3[216]=8'hab;
        mem_3[217]=8'ha9;
        mem_3[218]=8'haf;
        mem_3[219]=8'had;
        mem_3[220]=8'ha3;
        mem_3[221]=8'ha1;
        mem_3[222]=8'ha7;
        mem_3[223]=8'ha5;
        mem_3[224]=8'hdb;
        mem_3[225]=8'hd9;
        mem_3[226]=8'hdf;
        mem_3[227]=8'hdd;
        mem_3[228]=8'hd3;
        mem_3[229]=8'hd1;
        mem_3[230]=8'hd7;
        mem_3[231]=8'hd5;
        mem_3[232]=8'hcb;
        mem_3[233]=8'hc9;
        mem_3[234]=8'hcf;
        mem_3[235]=8'hcd;
        mem_3[236]=8'hc3;
        mem_3[237]=8'hc1;
        mem_3[238]=8'hc7;
        mem_3[239]=8'hc5;
        mem_3[240]=8'hfb;
        mem_3[241]=8'hf9;
        mem_3[242]=8'hff;
        mem_3[243]=8'hfd;
        mem_3[244]=8'hf3;
        mem_3[245]=8'hf1;
        mem_3[246]=8'hf7;
        mem_3[247]=8'hf5;
        mem_3[248]=8'heb;
        mem_3[249]=8'he9;
        mem_3[250]=8'hef;
        mem_3[251]=8'hed;
        mem_3[252]=8'he3;
        mem_3[253]=8'he1;
        mem_3[254]=8'he7;
        mem_3[255]=8'he5;
    end

    initial begin
        mem_4[0]=8'h0;
        mem_4[1]=8'h3;
        mem_4[2]=8'h6;
        mem_4[3]=8'h5;
        mem_4[4]=8'hc;
        mem_4[5]=8'hf;
        mem_4[6]=8'ha;
        mem_4[7]=8'h9;
        mem_4[8]=8'h18;
        mem_4[9]=8'h1b;
        mem_4[10]=8'h1e;
        mem_4[11]=8'h1d;
        mem_4[12]=8'h14;
        mem_4[13]=8'h17;
        mem_4[14]=8'h12;
        mem_4[15]=8'h11;
        mem_4[16]=8'h30;
        mem_4[17]=8'h33;
        mem_4[18]=8'h36;
        mem_4[19]=8'h35;
        mem_4[20]=8'h3c;
        mem_4[21]=8'h3f;
        mem_4[22]=8'h3a;
        mem_4[23]=8'h39;
        mem_4[24]=8'h28;
        mem_4[25]=8'h2b;
        mem_4[26]=8'h2e;
        mem_4[27]=8'h2d;
        mem_4[28]=8'h24;
        mem_4[29]=8'h27;
        mem_4[30]=8'h22;
        mem_4[31]=8'h21;
        mem_4[32]=8'h60;
        mem_4[33]=8'h63;
        mem_4[34]=8'h66;
        mem_4[35]=8'h65;
        mem_4[36]=8'h6c;
        mem_4[37]=8'h6f;
        mem_4[38]=8'h6a;
        mem_4[39]=8'h69;
        mem_4[40]=8'h78;
        mem_4[41]=8'h7b;
        mem_4[42]=8'h7e;
        mem_4[43]=8'h7d;
        mem_4[44]=8'h74;
        mem_4[45]=8'h77;
        mem_4[46]=8'h72;
        mem_4[47]=8'h71;
        mem_4[48]=8'h50;
        mem_4[49]=8'h53;
        mem_4[50]=8'h56;
        mem_4[51]=8'h55;
        mem_4[52]=8'h5c;
        mem_4[53]=8'h5f;
        mem_4[54]=8'h5a;
        mem_4[55]=8'h59;
        mem_4[56]=8'h48;
        mem_4[57]=8'h4b;
        mem_4[58]=8'h4e;
        mem_4[59]=8'h4d;
        mem_4[60]=8'h44;
        mem_4[61]=8'h47;
        mem_4[62]=8'h42;
        mem_4[63]=8'h41;
        mem_4[64]=8'hc0;
        mem_4[65]=8'hc3;
        mem_4[66]=8'hc6;
        mem_4[67]=8'hc5;
        mem_4[68]=8'hcc;
        mem_4[69]=8'hcf;
        mem_4[70]=8'hca;
        mem_4[71]=8'hc9;
        mem_4[72]=8'hd8;
        mem_4[73]=8'hdb;
        mem_4[74]=8'hde;
        mem_4[75]=8'hdd;
        mem_4[76]=8'hd4;
        mem_4[77]=8'hd7;
        mem_4[78]=8'hd2;
        mem_4[79]=8'hd1;
        mem_4[80]=8'hf0;
        mem_4[81]=8'hf3;
        mem_4[82]=8'hf6;
        mem_4[83]=8'hf5;
        mem_4[84]=8'hfc;
        mem_4[85]=8'hff;
        mem_4[86]=8'hfa;
        mem_4[87]=8'hf9;
        mem_4[88]=8'he8;
        mem_4[89]=8'heb;
        mem_4[90]=8'hee;
        mem_4[91]=8'hed;
        mem_4[92]=8'he4;
        mem_4[93]=8'he7;
        mem_4[94]=8'he2;
        mem_4[95]=8'he1;
        mem_4[96]=8'ha0;
        mem_4[97]=8'ha3;
        mem_4[98]=8'ha6;
        mem_4[99]=8'ha5;
        mem_4[100]=8'hac;
        mem_4[101]=8'haf;
        mem_4[102]=8'haa;
        mem_4[103]=8'ha9;
        mem_4[104]=8'hb8;
        mem_4[105]=8'hbb;
        mem_4[106]=8'hbe;
        mem_4[107]=8'hbd;
        mem_4[108]=8'hb4;
        mem_4[109]=8'hb7;
        mem_4[110]=8'hb2;
        mem_4[111]=8'hb1;
        mem_4[112]=8'h90;
        mem_4[113]=8'h93;
        mem_4[114]=8'h96;
        mem_4[115]=8'h95;
        mem_4[116]=8'h9c;
        mem_4[117]=8'h9f;
        mem_4[118]=8'h9a;
        mem_4[119]=8'h99;
        mem_4[120]=8'h88;
        mem_4[121]=8'h8b;
        mem_4[122]=8'h8e;
        mem_4[123]=8'h8d;
        mem_4[124]=8'h84;
        mem_4[125]=8'h87;
        mem_4[126]=8'h82;
        mem_4[127]=8'h81;
        mem_4[128]=8'h9b;
        mem_4[129]=8'h98;
        mem_4[130]=8'h9d;
        mem_4[131]=8'h9e;
        mem_4[132]=8'h97;
        mem_4[133]=8'h94;
        mem_4[134]=8'h91;
        mem_4[135]=8'h92;
        mem_4[136]=8'h83;
        mem_4[137]=8'h80;
        mem_4[138]=8'h85;
        mem_4[139]=8'h86;
        mem_4[140]=8'h8f;
        mem_4[141]=8'h8c;
        mem_4[142]=8'h89;
        mem_4[143]=8'h8a;
        mem_4[144]=8'hab;
        mem_4[145]=8'ha8;
        mem_4[146]=8'had;
        mem_4[147]=8'hae;
        mem_4[148]=8'ha7;
        mem_4[149]=8'ha4;
        mem_4[150]=8'ha1;
        mem_4[151]=8'ha2;
        mem_4[152]=8'hb3;
        mem_4[153]=8'hb0;
        mem_4[154]=8'hb5;
        mem_4[155]=8'hb6;
        mem_4[156]=8'hbf;
        mem_4[157]=8'hbc;
        mem_4[158]=8'hb9;
        mem_4[159]=8'hba;
        mem_4[160]=8'hfb;
        mem_4[161]=8'hf8;
        mem_4[162]=8'hfd;
        mem_4[163]=8'hfe;
        mem_4[164]=8'hf7;
        mem_4[165]=8'hf4;
        mem_4[166]=8'hf1;
        mem_4[167]=8'hf2;
        mem_4[168]=8'he3;
        mem_4[169]=8'he0;
        mem_4[170]=8'he5;
        mem_4[171]=8'he6;
        mem_4[172]=8'hef;
        mem_4[173]=8'hec;
        mem_4[174]=8'he9;
        mem_4[175]=8'hea;
        mem_4[176]=8'hcb;
        mem_4[177]=8'hc8;
        mem_4[178]=8'hcd;
        mem_4[179]=8'hce;
        mem_4[180]=8'hc7;
        mem_4[181]=8'hc4;
        mem_4[182]=8'hc1;
        mem_4[183]=8'hc2;
        mem_4[184]=8'hd3;
        mem_4[185]=8'hd0;
        mem_4[186]=8'hd5;
        mem_4[187]=8'hd6;
        mem_4[188]=8'hdf;
        mem_4[189]=8'hdc;
        mem_4[190]=8'hd9;
        mem_4[191]=8'hda;
        mem_4[192]=8'h5b;
        mem_4[193]=8'h58;
        mem_4[194]=8'h5d;
        mem_4[195]=8'h5e;
        mem_4[196]=8'h57;
        mem_4[197]=8'h54;
        mem_4[198]=8'h51;
        mem_4[199]=8'h52;
        mem_4[200]=8'h43;
        mem_4[201]=8'h40;
        mem_4[202]=8'h45;
        mem_4[203]=8'h46;
        mem_4[204]=8'h4f;
        mem_4[205]=8'h4c;
        mem_4[206]=8'h49;
        mem_4[207]=8'h4a;
        mem_4[208]=8'h6b;
        mem_4[209]=8'h68;
        mem_4[210]=8'h6d;
        mem_4[211]=8'h6e;
        mem_4[212]=8'h67;
        mem_4[213]=8'h64;
        mem_4[214]=8'h61;
        mem_4[215]=8'h62;
        mem_4[216]=8'h73;
        mem_4[217]=8'h70;
        mem_4[218]=8'h75;
        mem_4[219]=8'h76;
        mem_4[220]=8'h7f;
        mem_4[221]=8'h7c;
        mem_4[222]=8'h79;
        mem_4[223]=8'h7a;
        mem_4[224]=8'h3b;
        mem_4[225]=8'h38;
        mem_4[226]=8'h3d;
        mem_4[227]=8'h3e;
        mem_4[228]=8'h37;
        mem_4[229]=8'h34;
        mem_4[230]=8'h31;
        mem_4[231]=8'h32;
        mem_4[232]=8'h23;
        mem_4[233]=8'h20;
        mem_4[234]=8'h25;
        mem_4[235]=8'h26;
        mem_4[236]=8'h2f;
        mem_4[237]=8'h2c;
        mem_4[238]=8'h29;
        mem_4[239]=8'h2a;
        mem_4[240]=8'hb;
        mem_4[241]=8'h8;
        mem_4[242]=8'hd;
        mem_4[243]=8'he;
        mem_4[244]=8'h7;
        mem_4[245]=8'h4;
        mem_4[246]=8'h1;
        mem_4[247]=8'h2;
        mem_4[248]=8'h13;
        mem_4[249]=8'h10;
        mem_4[250]=8'h15;
        mem_4[251]=8'h16;
        mem_4[252]=8'h1f;
        mem_4[253]=8'h1c;
        mem_4[254]=8'h19;
        mem_4[255]=8'h1a;
    end

    initial begin
        mem_9[0]=8'h63;
        mem_9[1]=8'h7c;
        mem_9[2]=8'h77;
        mem_9[3]=8'h7b;
        mem_9[4]=8'hf2;
        mem_9[5]=8'h6b;
        mem_9[6]=8'h6f;
        mem_9[7]=8'hc5;
        mem_9[8]=8'h30;
        mem_9[9]=8'h1;
        mem_9[10]=8'h67;
        mem_9[11]=8'h2b;
        mem_9[12]=8'hfe;
        mem_9[13]=8'hd7;
        mem_9[14]=8'hab;
        mem_9[15]=8'h76;
        mem_9[16]=8'hca;
        mem_9[17]=8'h82;
        mem_9[18]=8'hc9;
        mem_9[19]=8'h7d;
        mem_9[20]=8'hfa;
        mem_9[21]=8'h59;
        mem_9[22]=8'h47;
        mem_9[23]=8'hf0;
        mem_9[24]=8'had;
        mem_9[25]=8'hd4;
        mem_9[26]=8'ha2;
        mem_9[27]=8'haf;
        mem_9[28]=8'h9c;
        mem_9[29]=8'ha4;
        mem_9[30]=8'h72;
        mem_9[31]=8'hc0;
        mem_9[32]=8'hb7;
        mem_9[33]=8'hfd;
        mem_9[34]=8'h93;
        mem_9[35]=8'h26;
        mem_9[36]=8'h36;
        mem_9[37]=8'h3f;
        mem_9[38]=8'hf7;
        mem_9[39]=8'hcc;
        mem_9[40]=8'h34;
        mem_9[41]=8'ha5;
        mem_9[42]=8'he5;
        mem_9[43]=8'hf1;
        mem_9[44]=8'h71;
        mem_9[45]=8'hd8;
        mem_9[46]=8'h31;
        mem_9[47]=8'h15;
        mem_9[48]=8'h4;
        mem_9[49]=8'hc7;
        mem_9[50]=8'h23;
        mem_9[51]=8'hc3;
        mem_9[52]=8'h18;
        mem_9[53]=8'h96;
        mem_9[54]=8'h5;
        mem_9[55]=8'h9a;
        mem_9[56]=8'h7;
        mem_9[57]=8'h12;
        mem_9[58]=8'h80;
        mem_9[59]=8'he2;
        mem_9[60]=8'heb;
        mem_9[61]=8'h27;
        mem_9[62]=8'hb2;
        mem_9[63]=8'h75;
        mem_9[64]=8'h9;
        mem_9[65]=8'h83;
        mem_9[66]=8'h2c;
        mem_9[67]=8'h1a;
        mem_9[68]=8'h1b;
        mem_9[69]=8'h6e;
        mem_9[70]=8'h5a;
        mem_9[71]=8'ha0;
        mem_9[72]=8'h52;
        mem_9[73]=8'h3b;
        mem_9[74]=8'hd6;
        mem_9[75]=8'hb3;
        mem_9[76]=8'h29;
        mem_9[77]=8'he3;
        mem_9[78]=8'h2f;
        mem_9[79]=8'h84;
        mem_9[80]=8'h53;
        mem_9[81]=8'hd1;
        mem_9[82]=8'h0;
        mem_9[83]=8'hed;
        mem_9[84]=8'h20;
        mem_9[85]=8'hfc;
        mem_9[86]=8'hb1;
        mem_9[87]=8'h5b;
        mem_9[88]=8'h6a;
        mem_9[89]=8'hcb;
        mem_9[90]=8'hbe;
        mem_9[91]=8'h39;
        mem_9[92]=8'h4a;
        mem_9[93]=8'h4c;
        mem_9[94]=8'h58;
        mem_9[95]=8'hcf;
        mem_9[96]=8'hd0;
        mem_9[97]=8'hef;
        mem_9[98]=8'haa;
        mem_9[99]=8'hfb;
        mem_9[100]=8'h43;
        mem_9[101]=8'h4d;
        mem_9[102]=8'h33;
        mem_9[103]=8'h85;
        mem_9[104]=8'h45;
        mem_9[105]=8'hf9;
        mem_9[106]=8'h2;
        mem_9[107]=8'h7f;
        mem_9[108]=8'h50;
        mem_9[109]=8'h3c;
        mem_9[110]=8'h9f;
        mem_9[111]=8'ha8;
        mem_9[112]=8'h51;
        mem_9[113]=8'ha3;
        mem_9[114]=8'h40;
        mem_9[115]=8'h8f;
        mem_9[116]=8'h92;
        mem_9[117]=8'h9d;
        mem_9[118]=8'h38;
        mem_9[119]=8'hf5;
        mem_9[120]=8'hbc;
        mem_9[121]=8'hb6;
        mem_9[122]=8'hda;
        mem_9[123]=8'h21;
        mem_9[124]=8'h10;
        mem_9[125]=8'hff;
        mem_9[126]=8'hf3;
        mem_9[127]=8'hd2;
        mem_9[128]=8'hcd;
        mem_9[129]=8'hc;
        mem_9[130]=8'h13;
        mem_9[131]=8'hec;
        mem_9[132]=8'h5f;
        mem_9[133]=8'h97;
        mem_9[134]=8'h44;
        mem_9[135]=8'h17;
        mem_9[136]=8'hc4;
        mem_9[137]=8'ha7;
        mem_9[138]=8'h7e;
        mem_9[139]=8'h3d;
        mem_9[140]=8'h64;
        mem_9[141]=8'h5d;
        mem_9[142]=8'h19;
        mem_9[143]=8'h73;
        mem_9[144]=8'h60;
        mem_9[145]=8'h81;
        mem_9[146]=8'h4f;
        mem_9[147]=8'hdc;
        mem_9[148]=8'h22;
        mem_9[149]=8'h2a;
        mem_9[150]=8'h90;
        mem_9[151]=8'h88;
        mem_9[152]=8'h46;
        mem_9[153]=8'hee;
        mem_9[154]=8'hb8;
        mem_9[155]=8'h14;
        mem_9[156]=8'hde;
        mem_9[157]=8'h5e;
        mem_9[158]=8'hb;
        mem_9[159]=8'hdb;
        mem_9[160]=8'he0;
        mem_9[161]=8'h32;
        mem_9[162]=8'h3a;
        mem_9[163]=8'ha;
        mem_9[164]=8'h49;
        mem_9[165]=8'h6;
        mem_9[166]=8'h24;
        mem_9[167]=8'h5c;
        mem_9[168]=8'hc2;
        mem_9[169]=8'hd3;
        mem_9[170]=8'hac;
        mem_9[171]=8'h62;
        mem_9[172]=8'h91;
        mem_9[173]=8'h95;
        mem_9[174]=8'he4;
        mem_9[175]=8'h79;
        mem_9[176]=8'he7;
        mem_9[177]=8'hc8;
        mem_9[178]=8'h37;
        mem_9[179]=8'h6d;
        mem_9[180]=8'h8d;
        mem_9[181]=8'hd5;
        mem_9[182]=8'h4e;
        mem_9[183]=8'ha9;
        mem_9[184]=8'h6c;
        mem_9[185]=8'h56;
        mem_9[186]=8'hf4;
        mem_9[187]=8'hea;
        mem_9[188]=8'h65;
        mem_9[189]=8'h7a;
        mem_9[190]=8'hae;
        mem_9[191]=8'h8;
        mem_9[192]=8'hba;
        mem_9[193]=8'h78;
        mem_9[194]=8'h25;
        mem_9[195]=8'h2e;
        mem_9[196]=8'h1c;
        mem_9[197]=8'ha6;
        mem_9[198]=8'hb4;
        mem_9[199]=8'hc6;
        mem_9[200]=8'he8;
        mem_9[201]=8'hdd;
        mem_9[202]=8'h74;
        mem_9[203]=8'h1f;
        mem_9[204]=8'h4b;
        mem_9[205]=8'hbd;
        mem_9[206]=8'h8b;
        mem_9[207]=8'h8a;
        mem_9[208]=8'h70;
        mem_9[209]=8'h3e;
        mem_9[210]=8'hb5;
        mem_9[211]=8'h66;
        mem_9[212]=8'h48;
        mem_9[213]=8'h3;
        mem_9[214]=8'hf6;
        mem_9[215]=8'he;
        mem_9[216]=8'h61;
        mem_9[217]=8'h35;
        mem_9[218]=8'h57;
        mem_9[219]=8'hb9;
        mem_9[220]=8'h86;
        mem_9[221]=8'hc1;
        mem_9[222]=8'h1d;
        mem_9[223]=8'h9e;
        mem_9[224]=8'he1;
        mem_9[225]=8'hf8;
        mem_9[226]=8'h98;
        mem_9[227]=8'h11;
        mem_9[228]=8'h69;
        mem_9[229]=8'hd9;
        mem_9[230]=8'h8e;
        mem_9[231]=8'h94;
        mem_9[232]=8'h9b;
        mem_9[233]=8'h1e;
        mem_9[234]=8'h87;
        mem_9[235]=8'he9;
        mem_9[236]=8'hce;
        mem_9[237]=8'h55;
        mem_9[238]=8'h28;
        mem_9[239]=8'hdf;
        mem_9[240]=8'h8c;
        mem_9[241]=8'ha1;
        mem_9[242]=8'h89;
        mem_9[243]=8'hd;
        mem_9[244]=8'hbf;
        mem_9[245]=8'he6;
        mem_9[246]=8'h42;
        mem_9[247]=8'h68;
        mem_9[248]=8'h41;
        mem_9[249]=8'h99;
        mem_9[250]=8'h2d;
        mem_9[251]=8'hf;
        mem_9[252]=8'hb0;
        mem_9[253]=8'h54;
        mem_9[254]=8'hbb;
        mem_9[255]=8'h16;
    end

    initial begin
        mem_10[0]=8'h63;
        mem_10[1]=8'h7c;
        mem_10[2]=8'h77;
        mem_10[3]=8'h7b;
        mem_10[4]=8'hf2;
        mem_10[5]=8'h6b;
        mem_10[6]=8'h6f;
        mem_10[7]=8'hc5;
        mem_10[8]=8'h30;
        mem_10[9]=8'h1;
        mem_10[10]=8'h67;
        mem_10[11]=8'h2b;
        mem_10[12]=8'hfe;
        mem_10[13]=8'hd7;
        mem_10[14]=8'hab;
        mem_10[15]=8'h76;
        mem_10[16]=8'hca;
        mem_10[17]=8'h82;
        mem_10[18]=8'hc9;
        mem_10[19]=8'h7d;
        mem_10[20]=8'hfa;
        mem_10[21]=8'h59;
        mem_10[22]=8'h47;
        mem_10[23]=8'hf0;
        mem_10[24]=8'had;
        mem_10[25]=8'hd4;
        mem_10[26]=8'ha2;
        mem_10[27]=8'haf;
        mem_10[28]=8'h9c;
        mem_10[29]=8'ha4;
        mem_10[30]=8'h72;
        mem_10[31]=8'hc0;
        mem_10[32]=8'hb7;
        mem_10[33]=8'hfd;
        mem_10[34]=8'h93;
        mem_10[35]=8'h26;
        mem_10[36]=8'h36;
        mem_10[37]=8'h3f;
        mem_10[38]=8'hf7;
        mem_10[39]=8'hcc;
        mem_10[40]=8'h34;
        mem_10[41]=8'ha5;
        mem_10[42]=8'he5;
        mem_10[43]=8'hf1;
        mem_10[44]=8'h71;
        mem_10[45]=8'hd8;
        mem_10[46]=8'h31;
        mem_10[47]=8'h15;
        mem_10[48]=8'h4;
        mem_10[49]=8'hc7;
        mem_10[50]=8'h23;
        mem_10[51]=8'hc3;
        mem_10[52]=8'h18;
        mem_10[53]=8'h96;
        mem_10[54]=8'h5;
        mem_10[55]=8'h9a;
        mem_10[56]=8'h7;
        mem_10[57]=8'h12;
        mem_10[58]=8'h80;
        mem_10[59]=8'he2;
        mem_10[60]=8'heb;
        mem_10[61]=8'h27;
        mem_10[62]=8'hb2;
        mem_10[63]=8'h75;
        mem_10[64]=8'h9;
        mem_10[65]=8'h83;
        mem_10[66]=8'h2c;
        mem_10[67]=8'h1a;
        mem_10[68]=8'h1b;
        mem_10[69]=8'h6e;
        mem_10[70]=8'h5a;
        mem_10[71]=8'ha0;
        mem_10[72]=8'h52;
        mem_10[73]=8'h3b;
        mem_10[74]=8'hd6;
        mem_10[75]=8'hb3;
        mem_10[76]=8'h29;
        mem_10[77]=8'he3;
        mem_10[78]=8'h2f;
        mem_10[79]=8'h84;
        mem_10[80]=8'h53;
        mem_10[81]=8'hd1;
        mem_10[82]=8'h0;
        mem_10[83]=8'hed;
        mem_10[84]=8'h20;
        mem_10[85]=8'hfc;
        mem_10[86]=8'hb1;
        mem_10[87]=8'h5b;
        mem_10[88]=8'h6a;
        mem_10[89]=8'hcb;
        mem_10[90]=8'hbe;
        mem_10[91]=8'h39;
        mem_10[92]=8'h4a;
        mem_10[93]=8'h4c;
        mem_10[94]=8'h58;
        mem_10[95]=8'hcf;
        mem_10[96]=8'hd0;
        mem_10[97]=8'hef;
        mem_10[98]=8'haa;
        mem_10[99]=8'hfb;
        mem_10[100]=8'h43;
        mem_10[101]=8'h4d;
        mem_10[102]=8'h33;
        mem_10[103]=8'h85;
        mem_10[104]=8'h45;
        mem_10[105]=8'hf9;
        mem_10[106]=8'h2;
        mem_10[107]=8'h7f;
        mem_10[108]=8'h50;
        mem_10[109]=8'h3c;
        mem_10[110]=8'h9f;
        mem_10[111]=8'ha8;
        mem_10[112]=8'h51;
        mem_10[113]=8'ha3;
        mem_10[114]=8'h40;
        mem_10[115]=8'h8f;
        mem_10[116]=8'h92;
        mem_10[117]=8'h9d;
        mem_10[118]=8'h38;
        mem_10[119]=8'hf5;
        mem_10[120]=8'hbc;
        mem_10[121]=8'hb6;
        mem_10[122]=8'hda;
        mem_10[123]=8'h21;
        mem_10[124]=8'h10;
        mem_10[125]=8'hff;
        mem_10[126]=8'hf3;
        mem_10[127]=8'hd2;
        mem_10[128]=8'hcd;
        mem_10[129]=8'hc;
        mem_10[130]=8'h13;
        mem_10[131]=8'hec;
        mem_10[132]=8'h5f;
        mem_10[133]=8'h97;
        mem_10[134]=8'h44;
        mem_10[135]=8'h17;
        mem_10[136]=8'hc4;
        mem_10[137]=8'ha7;
        mem_10[138]=8'h7e;
        mem_10[139]=8'h3d;
        mem_10[140]=8'h64;
        mem_10[141]=8'h5d;
        mem_10[142]=8'h19;
        mem_10[143]=8'h73;
        mem_10[144]=8'h60;
        mem_10[145]=8'h81;
        mem_10[146]=8'h4f;
        mem_10[147]=8'hdc;
        mem_10[148]=8'h22;
        mem_10[149]=8'h2a;
        mem_10[150]=8'h90;
        mem_10[151]=8'h88;
        mem_10[152]=8'h46;
        mem_10[153]=8'hee;
        mem_10[154]=8'hb8;
        mem_10[155]=8'h14;
        mem_10[156]=8'hde;
        mem_10[157]=8'h5e;
        mem_10[158]=8'hb;
        mem_10[159]=8'hdb;
        mem_10[160]=8'he0;
        mem_10[161]=8'h32;
        mem_10[162]=8'h3a;
        mem_10[163]=8'ha;
        mem_10[164]=8'h49;
        mem_10[165]=8'h6;
        mem_10[166]=8'h24;
        mem_10[167]=8'h5c;
        mem_10[168]=8'hc2;
        mem_10[169]=8'hd3;
        mem_10[170]=8'hac;
        mem_10[171]=8'h62;
        mem_10[172]=8'h91;
        mem_10[173]=8'h95;
        mem_10[174]=8'he4;
        mem_10[175]=8'h79;
        mem_10[176]=8'he7;
        mem_10[177]=8'hc8;
        mem_10[178]=8'h37;
        mem_10[179]=8'h6d;
        mem_10[180]=8'h8d;
        mem_10[181]=8'hd5;
        mem_10[182]=8'h4e;
        mem_10[183]=8'ha9;
        mem_10[184]=8'h6c;
        mem_10[185]=8'h56;
        mem_10[186]=8'hf4;
        mem_10[187]=8'hea;
        mem_10[188]=8'h65;
        mem_10[189]=8'h7a;
        mem_10[190]=8'hae;
        mem_10[191]=8'h8;
        mem_10[192]=8'hba;
        mem_10[193]=8'h78;
        mem_10[194]=8'h25;
        mem_10[195]=8'h2e;
        mem_10[196]=8'h1c;
        mem_10[197]=8'ha6;
        mem_10[198]=8'hb4;
        mem_10[199]=8'hc6;
        mem_10[200]=8'he8;
        mem_10[201]=8'hdd;
        mem_10[202]=8'h74;
        mem_10[203]=8'h1f;
        mem_10[204]=8'h4b;
        mem_10[205]=8'hbd;
        mem_10[206]=8'h8b;
        mem_10[207]=8'h8a;
        mem_10[208]=8'h70;
        mem_10[209]=8'h3e;
        mem_10[210]=8'hb5;
        mem_10[211]=8'h66;
        mem_10[212]=8'h48;
        mem_10[213]=8'h3;
        mem_10[214]=8'hf6;
        mem_10[215]=8'he;
        mem_10[216]=8'h61;
        mem_10[217]=8'h35;
        mem_10[218]=8'h57;
        mem_10[219]=8'hb9;
        mem_10[220]=8'h86;
        mem_10[221]=8'hc1;
        mem_10[222]=8'h1d;
        mem_10[223]=8'h9e;
        mem_10[224]=8'he1;
        mem_10[225]=8'hf8;
        mem_10[226]=8'h98;
        mem_10[227]=8'h11;
        mem_10[228]=8'h69;
        mem_10[229]=8'hd9;
        mem_10[230]=8'h8e;
        mem_10[231]=8'h94;
        mem_10[232]=8'h9b;
        mem_10[233]=8'h1e;
        mem_10[234]=8'h87;
        mem_10[235]=8'he9;
        mem_10[236]=8'hce;
        mem_10[237]=8'h55;
        mem_10[238]=8'h28;
        mem_10[239]=8'hdf;
        mem_10[240]=8'h8c;
        mem_10[241]=8'ha1;
        mem_10[242]=8'h89;
        mem_10[243]=8'hd;
        mem_10[244]=8'hbf;
        mem_10[245]=8'he6;
        mem_10[246]=8'h42;
        mem_10[247]=8'h68;
        mem_10[248]=8'h41;
        mem_10[249]=8'h99;
        mem_10[250]=8'h2d;
        mem_10[251]=8'hf;
        mem_10[252]=8'hb0;
        mem_10[253]=8'h54;
        mem_10[254]=8'hbb;
        mem_10[255]=8'h16;
    end

    initial begin
        mem_11[0]=8'h63;
        mem_11[1]=8'h7c;
        mem_11[2]=8'h77;
        mem_11[3]=8'h7b;
        mem_11[4]=8'hf2;
        mem_11[5]=8'h6b;
        mem_11[6]=8'h6f;
        mem_11[7]=8'hc5;
        mem_11[8]=8'h30;
        mem_11[9]=8'h1;
        mem_11[10]=8'h67;
        mem_11[11]=8'h2b;
        mem_11[12]=8'hfe;
        mem_11[13]=8'hd7;
        mem_11[14]=8'hab;
        mem_11[15]=8'h76;
        mem_11[16]=8'hca;
        mem_11[17]=8'h82;
        mem_11[18]=8'hc9;
        mem_11[19]=8'h7d;
        mem_11[20]=8'hfa;
        mem_11[21]=8'h59;
        mem_11[22]=8'h47;
        mem_11[23]=8'hf0;
        mem_11[24]=8'had;
        mem_11[25]=8'hd4;
        mem_11[26]=8'ha2;
        mem_11[27]=8'haf;
        mem_11[28]=8'h9c;
        mem_11[29]=8'ha4;
        mem_11[30]=8'h72;
        mem_11[31]=8'hc0;
        mem_11[32]=8'hb7;
        mem_11[33]=8'hfd;
        mem_11[34]=8'h93;
        mem_11[35]=8'h26;
        mem_11[36]=8'h36;
        mem_11[37]=8'h3f;
        mem_11[38]=8'hf7;
        mem_11[39]=8'hcc;
        mem_11[40]=8'h34;
        mem_11[41]=8'ha5;
        mem_11[42]=8'he5;
        mem_11[43]=8'hf1;
        mem_11[44]=8'h71;
        mem_11[45]=8'hd8;
        mem_11[46]=8'h31;
        mem_11[47]=8'h15;
        mem_11[48]=8'h4;
        mem_11[49]=8'hc7;
        mem_11[50]=8'h23;
        mem_11[51]=8'hc3;
        mem_11[52]=8'h18;
        mem_11[53]=8'h96;
        mem_11[54]=8'h5;
        mem_11[55]=8'h9a;
        mem_11[56]=8'h7;
        mem_11[57]=8'h12;
        mem_11[58]=8'h80;
        mem_11[59]=8'he2;
        mem_11[60]=8'heb;
        mem_11[61]=8'h27;
        mem_11[62]=8'hb2;
        mem_11[63]=8'h75;
        mem_11[64]=8'h9;
        mem_11[65]=8'h83;
        mem_11[66]=8'h2c;
        mem_11[67]=8'h1a;
        mem_11[68]=8'h1b;
        mem_11[69]=8'h6e;
        mem_11[70]=8'h5a;
        mem_11[71]=8'ha0;
        mem_11[72]=8'h52;
        mem_11[73]=8'h3b;
        mem_11[74]=8'hd6;
        mem_11[75]=8'hb3;
        mem_11[76]=8'h29;
        mem_11[77]=8'he3;
        mem_11[78]=8'h2f;
        mem_11[79]=8'h84;
        mem_11[80]=8'h53;
        mem_11[81]=8'hd1;
        mem_11[82]=8'h0;
        mem_11[83]=8'hed;
        mem_11[84]=8'h20;
        mem_11[85]=8'hfc;
        mem_11[86]=8'hb1;
        mem_11[87]=8'h5b;
        mem_11[88]=8'h6a;
        mem_11[89]=8'hcb;
        mem_11[90]=8'hbe;
        mem_11[91]=8'h39;
        mem_11[92]=8'h4a;
        mem_11[93]=8'h4c;
        mem_11[94]=8'h58;
        mem_11[95]=8'hcf;
        mem_11[96]=8'hd0;
        mem_11[97]=8'hef;
        mem_11[98]=8'haa;
        mem_11[99]=8'hfb;
        mem_11[100]=8'h43;
        mem_11[101]=8'h4d;
        mem_11[102]=8'h33;
        mem_11[103]=8'h85;
        mem_11[104]=8'h45;
        mem_11[105]=8'hf9;
        mem_11[106]=8'h2;
        mem_11[107]=8'h7f;
        mem_11[108]=8'h50;
        mem_11[109]=8'h3c;
        mem_11[110]=8'h9f;
        mem_11[111]=8'ha8;
        mem_11[112]=8'h51;
        mem_11[113]=8'ha3;
        mem_11[114]=8'h40;
        mem_11[115]=8'h8f;
        mem_11[116]=8'h92;
        mem_11[117]=8'h9d;
        mem_11[118]=8'h38;
        mem_11[119]=8'hf5;
        mem_11[120]=8'hbc;
        mem_11[121]=8'hb6;
        mem_11[122]=8'hda;
        mem_11[123]=8'h21;
        mem_11[124]=8'h10;
        mem_11[125]=8'hff;
        mem_11[126]=8'hf3;
        mem_11[127]=8'hd2;
        mem_11[128]=8'hcd;
        mem_11[129]=8'hc;
        mem_11[130]=8'h13;
        mem_11[131]=8'hec;
        mem_11[132]=8'h5f;
        mem_11[133]=8'h97;
        mem_11[134]=8'h44;
        mem_11[135]=8'h17;
        mem_11[136]=8'hc4;
        mem_11[137]=8'ha7;
        mem_11[138]=8'h7e;
        mem_11[139]=8'h3d;
        mem_11[140]=8'h64;
        mem_11[141]=8'h5d;
        mem_11[142]=8'h19;
        mem_11[143]=8'h73;
        mem_11[144]=8'h60;
        mem_11[145]=8'h81;
        mem_11[146]=8'h4f;
        mem_11[147]=8'hdc;
        mem_11[148]=8'h22;
        mem_11[149]=8'h2a;
        mem_11[150]=8'h90;
        mem_11[151]=8'h88;
        mem_11[152]=8'h46;
        mem_11[153]=8'hee;
        mem_11[154]=8'hb8;
        mem_11[155]=8'h14;
        mem_11[156]=8'hde;
        mem_11[157]=8'h5e;
        mem_11[158]=8'hb;
        mem_11[159]=8'hdb;
        mem_11[160]=8'he0;
        mem_11[161]=8'h32;
        mem_11[162]=8'h3a;
        mem_11[163]=8'ha;
        mem_11[164]=8'h49;
        mem_11[165]=8'h6;
        mem_11[166]=8'h24;
        mem_11[167]=8'h5c;
        mem_11[168]=8'hc2;
        mem_11[169]=8'hd3;
        mem_11[170]=8'hac;
        mem_11[171]=8'h62;
        mem_11[172]=8'h91;
        mem_11[173]=8'h95;
        mem_11[174]=8'he4;
        mem_11[175]=8'h79;
        mem_11[176]=8'he7;
        mem_11[177]=8'hc8;
        mem_11[178]=8'h37;
        mem_11[179]=8'h6d;
        mem_11[180]=8'h8d;
        mem_11[181]=8'hd5;
        mem_11[182]=8'h4e;
        mem_11[183]=8'ha9;
        mem_11[184]=8'h6c;
        mem_11[185]=8'h56;
        mem_11[186]=8'hf4;
        mem_11[187]=8'hea;
        mem_11[188]=8'h65;
        mem_11[189]=8'h7a;
        mem_11[190]=8'hae;
        mem_11[191]=8'h8;
        mem_11[192]=8'hba;
        mem_11[193]=8'h78;
        mem_11[194]=8'h25;
        mem_11[195]=8'h2e;
        mem_11[196]=8'h1c;
        mem_11[197]=8'ha6;
        mem_11[198]=8'hb4;
        mem_11[199]=8'hc6;
        mem_11[200]=8'he8;
        mem_11[201]=8'hdd;
        mem_11[202]=8'h74;
        mem_11[203]=8'h1f;
        mem_11[204]=8'h4b;
        mem_11[205]=8'hbd;
        mem_11[206]=8'h8b;
        mem_11[207]=8'h8a;
        mem_11[208]=8'h70;
        mem_11[209]=8'h3e;
        mem_11[210]=8'hb5;
        mem_11[211]=8'h66;
        mem_11[212]=8'h48;
        mem_11[213]=8'h3;
        mem_11[214]=8'hf6;
        mem_11[215]=8'he;
        mem_11[216]=8'h61;
        mem_11[217]=8'h35;
        mem_11[218]=8'h57;
        mem_11[219]=8'hb9;
        mem_11[220]=8'h86;
        mem_11[221]=8'hc1;
        mem_11[222]=8'h1d;
        mem_11[223]=8'h9e;
        mem_11[224]=8'he1;
        mem_11[225]=8'hf8;
        mem_11[226]=8'h98;
        mem_11[227]=8'h11;
        mem_11[228]=8'h69;
        mem_11[229]=8'hd9;
        mem_11[230]=8'h8e;
        mem_11[231]=8'h94;
        mem_11[232]=8'h9b;
        mem_11[233]=8'h1e;
        mem_11[234]=8'h87;
        mem_11[235]=8'he9;
        mem_11[236]=8'hce;
        mem_11[237]=8'h55;
        mem_11[238]=8'h28;
        mem_11[239]=8'hdf;
        mem_11[240]=8'h8c;
        mem_11[241]=8'ha1;
        mem_11[242]=8'h89;
        mem_11[243]=8'hd;
        mem_11[244]=8'hbf;
        mem_11[245]=8'he6;
        mem_11[246]=8'h42;
        mem_11[247]=8'h68;
        mem_11[248]=8'h41;
        mem_11[249]=8'h99;
        mem_11[250]=8'h2d;
        mem_11[251]=8'hf;
        mem_11[252]=8'hb0;
        mem_11[253]=8'h54;
        mem_11[254]=8'hbb;
        mem_11[255]=8'h16;
    end

    initial begin
        mem_12[0]=8'h63;
        mem_12[1]=8'h7c;
        mem_12[2]=8'h77;
        mem_12[3]=8'h7b;
        mem_12[4]=8'hf2;
        mem_12[5]=8'h6b;
        mem_12[6]=8'h6f;
        mem_12[7]=8'hc5;
        mem_12[8]=8'h30;
        mem_12[9]=8'h1;
        mem_12[10]=8'h67;
        mem_12[11]=8'h2b;
        mem_12[12]=8'hfe;
        mem_12[13]=8'hd7;
        mem_12[14]=8'hab;
        mem_12[15]=8'h76;
        mem_12[16]=8'hca;
        mem_12[17]=8'h82;
        mem_12[18]=8'hc9;
        mem_12[19]=8'h7d;
        mem_12[20]=8'hfa;
        mem_12[21]=8'h59;
        mem_12[22]=8'h47;
        mem_12[23]=8'hf0;
        mem_12[24]=8'had;
        mem_12[25]=8'hd4;
        mem_12[26]=8'ha2;
        mem_12[27]=8'haf;
        mem_12[28]=8'h9c;
        mem_12[29]=8'ha4;
        mem_12[30]=8'h72;
        mem_12[31]=8'hc0;
        mem_12[32]=8'hb7;
        mem_12[33]=8'hfd;
        mem_12[34]=8'h93;
        mem_12[35]=8'h26;
        mem_12[36]=8'h36;
        mem_12[37]=8'h3f;
        mem_12[38]=8'hf7;
        mem_12[39]=8'hcc;
        mem_12[40]=8'h34;
        mem_12[41]=8'ha5;
        mem_12[42]=8'he5;
        mem_12[43]=8'hf1;
        mem_12[44]=8'h71;
        mem_12[45]=8'hd8;
        mem_12[46]=8'h31;
        mem_12[47]=8'h15;
        mem_12[48]=8'h4;
        mem_12[49]=8'hc7;
        mem_12[50]=8'h23;
        mem_12[51]=8'hc3;
        mem_12[52]=8'h18;
        mem_12[53]=8'h96;
        mem_12[54]=8'h5;
        mem_12[55]=8'h9a;
        mem_12[56]=8'h7;
        mem_12[57]=8'h12;
        mem_12[58]=8'h80;
        mem_12[59]=8'he2;
        mem_12[60]=8'heb;
        mem_12[61]=8'h27;
        mem_12[62]=8'hb2;
        mem_12[63]=8'h75;
        mem_12[64]=8'h9;
        mem_12[65]=8'h83;
        mem_12[66]=8'h2c;
        mem_12[67]=8'h1a;
        mem_12[68]=8'h1b;
        mem_12[69]=8'h6e;
        mem_12[70]=8'h5a;
        mem_12[71]=8'ha0;
        mem_12[72]=8'h52;
        mem_12[73]=8'h3b;
        mem_12[74]=8'hd6;
        mem_12[75]=8'hb3;
        mem_12[76]=8'h29;
        mem_12[77]=8'he3;
        mem_12[78]=8'h2f;
        mem_12[79]=8'h84;
        mem_12[80]=8'h53;
        mem_12[81]=8'hd1;
        mem_12[82]=8'h0;
        mem_12[83]=8'hed;
        mem_12[84]=8'h20;
        mem_12[85]=8'hfc;
        mem_12[86]=8'hb1;
        mem_12[87]=8'h5b;
        mem_12[88]=8'h6a;
        mem_12[89]=8'hcb;
        mem_12[90]=8'hbe;
        mem_12[91]=8'h39;
        mem_12[92]=8'h4a;
        mem_12[93]=8'h4c;
        mem_12[94]=8'h58;
        mem_12[95]=8'hcf;
        mem_12[96]=8'hd0;
        mem_12[97]=8'hef;
        mem_12[98]=8'haa;
        mem_12[99]=8'hfb;
        mem_12[100]=8'h43;
        mem_12[101]=8'h4d;
        mem_12[102]=8'h33;
        mem_12[103]=8'h85;
        mem_12[104]=8'h45;
        mem_12[105]=8'hf9;
        mem_12[106]=8'h2;
        mem_12[107]=8'h7f;
        mem_12[108]=8'h50;
        mem_12[109]=8'h3c;
        mem_12[110]=8'h9f;
        mem_12[111]=8'ha8;
        mem_12[112]=8'h51;
        mem_12[113]=8'ha3;
        mem_12[114]=8'h40;
        mem_12[115]=8'h8f;
        mem_12[116]=8'h92;
        mem_12[117]=8'h9d;
        mem_12[118]=8'h38;
        mem_12[119]=8'hf5;
        mem_12[120]=8'hbc;
        mem_12[121]=8'hb6;
        mem_12[122]=8'hda;
        mem_12[123]=8'h21;
        mem_12[124]=8'h10;
        mem_12[125]=8'hff;
        mem_12[126]=8'hf3;
        mem_12[127]=8'hd2;
        mem_12[128]=8'hcd;
        mem_12[129]=8'hc;
        mem_12[130]=8'h13;
        mem_12[131]=8'hec;
        mem_12[132]=8'h5f;
        mem_12[133]=8'h97;
        mem_12[134]=8'h44;
        mem_12[135]=8'h17;
        mem_12[136]=8'hc4;
        mem_12[137]=8'ha7;
        mem_12[138]=8'h7e;
        mem_12[139]=8'h3d;
        mem_12[140]=8'h64;
        mem_12[141]=8'h5d;
        mem_12[142]=8'h19;
        mem_12[143]=8'h73;
        mem_12[144]=8'h60;
        mem_12[145]=8'h81;
        mem_12[146]=8'h4f;
        mem_12[147]=8'hdc;
        mem_12[148]=8'h22;
        mem_12[149]=8'h2a;
        mem_12[150]=8'h90;
        mem_12[151]=8'h88;
        mem_12[152]=8'h46;
        mem_12[153]=8'hee;
        mem_12[154]=8'hb8;
        mem_12[155]=8'h14;
        mem_12[156]=8'hde;
        mem_12[157]=8'h5e;
        mem_12[158]=8'hb;
        mem_12[159]=8'hdb;
        mem_12[160]=8'he0;
        mem_12[161]=8'h32;
        mem_12[162]=8'h3a;
        mem_12[163]=8'ha;
        mem_12[164]=8'h49;
        mem_12[165]=8'h6;
        mem_12[166]=8'h24;
        mem_12[167]=8'h5c;
        mem_12[168]=8'hc2;
        mem_12[169]=8'hd3;
        mem_12[170]=8'hac;
        mem_12[171]=8'h62;
        mem_12[172]=8'h91;
        mem_12[173]=8'h95;
        mem_12[174]=8'he4;
        mem_12[175]=8'h79;
        mem_12[176]=8'he7;
        mem_12[177]=8'hc8;
        mem_12[178]=8'h37;
        mem_12[179]=8'h6d;
        mem_12[180]=8'h8d;
        mem_12[181]=8'hd5;
        mem_12[182]=8'h4e;
        mem_12[183]=8'ha9;
        mem_12[184]=8'h6c;
        mem_12[185]=8'h56;
        mem_12[186]=8'hf4;
        mem_12[187]=8'hea;
        mem_12[188]=8'h65;
        mem_12[189]=8'h7a;
        mem_12[190]=8'hae;
        mem_12[191]=8'h8;
        mem_12[192]=8'hba;
        mem_12[193]=8'h78;
        mem_12[194]=8'h25;
        mem_12[195]=8'h2e;
        mem_12[196]=8'h1c;
        mem_12[197]=8'ha6;
        mem_12[198]=8'hb4;
        mem_12[199]=8'hc6;
        mem_12[200]=8'he8;
        mem_12[201]=8'hdd;
        mem_12[202]=8'h74;
        mem_12[203]=8'h1f;
        mem_12[204]=8'h4b;
        mem_12[205]=8'hbd;
        mem_12[206]=8'h8b;
        mem_12[207]=8'h8a;
        mem_12[208]=8'h70;
        mem_12[209]=8'h3e;
        mem_12[210]=8'hb5;
        mem_12[211]=8'h66;
        mem_12[212]=8'h48;
        mem_12[213]=8'h3;
        mem_12[214]=8'hf6;
        mem_12[215]=8'he;
        mem_12[216]=8'h61;
        mem_12[217]=8'h35;
        mem_12[218]=8'h57;
        mem_12[219]=8'hb9;
        mem_12[220]=8'h86;
        mem_12[221]=8'hc1;
        mem_12[222]=8'h1d;
        mem_12[223]=8'h9e;
        mem_12[224]=8'he1;
        mem_12[225]=8'hf8;
        mem_12[226]=8'h98;
        mem_12[227]=8'h11;
        mem_12[228]=8'h69;
        mem_12[229]=8'hd9;
        mem_12[230]=8'h8e;
        mem_12[231]=8'h94;
        mem_12[232]=8'h9b;
        mem_12[233]=8'h1e;
        mem_12[234]=8'h87;
        mem_12[235]=8'he9;
        mem_12[236]=8'hce;
        mem_12[237]=8'h55;
        mem_12[238]=8'h28;
        mem_12[239]=8'hdf;
        mem_12[240]=8'h8c;
        mem_12[241]=8'ha1;
        mem_12[242]=8'h89;
        mem_12[243]=8'hd;
        mem_12[244]=8'hbf;
        mem_12[245]=8'he6;
        mem_12[246]=8'h42;
        mem_12[247]=8'h68;
        mem_12[248]=8'h41;
        mem_12[249]=8'h99;
        mem_12[250]=8'h2d;
        mem_12[251]=8'hf;
        mem_12[252]=8'hb0;
        mem_12[253]=8'h54;
        mem_12[254]=8'hbb;
        mem_12[255]=8'h16;
    end

    initial begin
        mem_13[0]=8'h63;
        mem_13[1]=8'h7c;
        mem_13[2]=8'h77;
        mem_13[3]=8'h7b;
        mem_13[4]=8'hf2;
        mem_13[5]=8'h6b;
        mem_13[6]=8'h6f;
        mem_13[7]=8'hc5;
        mem_13[8]=8'h30;
        mem_13[9]=8'h1;
        mem_13[10]=8'h67;
        mem_13[11]=8'h2b;
        mem_13[12]=8'hfe;
        mem_13[13]=8'hd7;
        mem_13[14]=8'hab;
        mem_13[15]=8'h76;
        mem_13[16]=8'hca;
        mem_13[17]=8'h82;
        mem_13[18]=8'hc9;
        mem_13[19]=8'h7d;
        mem_13[20]=8'hfa;
        mem_13[21]=8'h59;
        mem_13[22]=8'h47;
        mem_13[23]=8'hf0;
        mem_13[24]=8'had;
        mem_13[25]=8'hd4;
        mem_13[26]=8'ha2;
        mem_13[27]=8'haf;
        mem_13[28]=8'h9c;
        mem_13[29]=8'ha4;
        mem_13[30]=8'h72;
        mem_13[31]=8'hc0;
        mem_13[32]=8'hb7;
        mem_13[33]=8'hfd;
        mem_13[34]=8'h93;
        mem_13[35]=8'h26;
        mem_13[36]=8'h36;
        mem_13[37]=8'h3f;
        mem_13[38]=8'hf7;
        mem_13[39]=8'hcc;
        mem_13[40]=8'h34;
        mem_13[41]=8'ha5;
        mem_13[42]=8'he5;
        mem_13[43]=8'hf1;
        mem_13[44]=8'h71;
        mem_13[45]=8'hd8;
        mem_13[46]=8'h31;
        mem_13[47]=8'h15;
        mem_13[48]=8'h4;
        mem_13[49]=8'hc7;
        mem_13[50]=8'h23;
        mem_13[51]=8'hc3;
        mem_13[52]=8'h18;
        mem_13[53]=8'h96;
        mem_13[54]=8'h5;
        mem_13[55]=8'h9a;
        mem_13[56]=8'h7;
        mem_13[57]=8'h12;
        mem_13[58]=8'h80;
        mem_13[59]=8'he2;
        mem_13[60]=8'heb;
        mem_13[61]=8'h27;
        mem_13[62]=8'hb2;
        mem_13[63]=8'h75;
        mem_13[64]=8'h9;
        mem_13[65]=8'h83;
        mem_13[66]=8'h2c;
        mem_13[67]=8'h1a;
        mem_13[68]=8'h1b;
        mem_13[69]=8'h6e;
        mem_13[70]=8'h5a;
        mem_13[71]=8'ha0;
        mem_13[72]=8'h52;
        mem_13[73]=8'h3b;
        mem_13[74]=8'hd6;
        mem_13[75]=8'hb3;
        mem_13[76]=8'h29;
        mem_13[77]=8'he3;
        mem_13[78]=8'h2f;
        mem_13[79]=8'h84;
        mem_13[80]=8'h53;
        mem_13[81]=8'hd1;
        mem_13[82]=8'h0;
        mem_13[83]=8'hed;
        mem_13[84]=8'h20;
        mem_13[85]=8'hfc;
        mem_13[86]=8'hb1;
        mem_13[87]=8'h5b;
        mem_13[88]=8'h6a;
        mem_13[89]=8'hcb;
        mem_13[90]=8'hbe;
        mem_13[91]=8'h39;
        mem_13[92]=8'h4a;
        mem_13[93]=8'h4c;
        mem_13[94]=8'h58;
        mem_13[95]=8'hcf;
        mem_13[96]=8'hd0;
        mem_13[97]=8'hef;
        mem_13[98]=8'haa;
        mem_13[99]=8'hfb;
        mem_13[100]=8'h43;
        mem_13[101]=8'h4d;
        mem_13[102]=8'h33;
        mem_13[103]=8'h85;
        mem_13[104]=8'h45;
        mem_13[105]=8'hf9;
        mem_13[106]=8'h2;
        mem_13[107]=8'h7f;
        mem_13[108]=8'h50;
        mem_13[109]=8'h3c;
        mem_13[110]=8'h9f;
        mem_13[111]=8'ha8;
        mem_13[112]=8'h51;
        mem_13[113]=8'ha3;
        mem_13[114]=8'h40;
        mem_13[115]=8'h8f;
        mem_13[116]=8'h92;
        mem_13[117]=8'h9d;
        mem_13[118]=8'h38;
        mem_13[119]=8'hf5;
        mem_13[120]=8'hbc;
        mem_13[121]=8'hb6;
        mem_13[122]=8'hda;
        mem_13[123]=8'h21;
        mem_13[124]=8'h10;
        mem_13[125]=8'hff;
        mem_13[126]=8'hf3;
        mem_13[127]=8'hd2;
        mem_13[128]=8'hcd;
        mem_13[129]=8'hc;
        mem_13[130]=8'h13;
        mem_13[131]=8'hec;
        mem_13[132]=8'h5f;
        mem_13[133]=8'h97;
        mem_13[134]=8'h44;
        mem_13[135]=8'h17;
        mem_13[136]=8'hc4;
        mem_13[137]=8'ha7;
        mem_13[138]=8'h7e;
        mem_13[139]=8'h3d;
        mem_13[140]=8'h64;
        mem_13[141]=8'h5d;
        mem_13[142]=8'h19;
        mem_13[143]=8'h73;
        mem_13[144]=8'h60;
        mem_13[145]=8'h81;
        mem_13[146]=8'h4f;
        mem_13[147]=8'hdc;
        mem_13[148]=8'h22;
        mem_13[149]=8'h2a;
        mem_13[150]=8'h90;
        mem_13[151]=8'h88;
        mem_13[152]=8'h46;
        mem_13[153]=8'hee;
        mem_13[154]=8'hb8;
        mem_13[155]=8'h14;
        mem_13[156]=8'hde;
        mem_13[157]=8'h5e;
        mem_13[158]=8'hb;
        mem_13[159]=8'hdb;
        mem_13[160]=8'he0;
        mem_13[161]=8'h32;
        mem_13[162]=8'h3a;
        mem_13[163]=8'ha;
        mem_13[164]=8'h49;
        mem_13[165]=8'h6;
        mem_13[166]=8'h24;
        mem_13[167]=8'h5c;
        mem_13[168]=8'hc2;
        mem_13[169]=8'hd3;
        mem_13[170]=8'hac;
        mem_13[171]=8'h62;
        mem_13[172]=8'h91;
        mem_13[173]=8'h95;
        mem_13[174]=8'he4;
        mem_13[175]=8'h79;
        mem_13[176]=8'he7;
        mem_13[177]=8'hc8;
        mem_13[178]=8'h37;
        mem_13[179]=8'h6d;
        mem_13[180]=8'h8d;
        mem_13[181]=8'hd5;
        mem_13[182]=8'h4e;
        mem_13[183]=8'ha9;
        mem_13[184]=8'h6c;
        mem_13[185]=8'h56;
        mem_13[186]=8'hf4;
        mem_13[187]=8'hea;
        mem_13[188]=8'h65;
        mem_13[189]=8'h7a;
        mem_13[190]=8'hae;
        mem_13[191]=8'h8;
        mem_13[192]=8'hba;
        mem_13[193]=8'h78;
        mem_13[194]=8'h25;
        mem_13[195]=8'h2e;
        mem_13[196]=8'h1c;
        mem_13[197]=8'ha6;
        mem_13[198]=8'hb4;
        mem_13[199]=8'hc6;
        mem_13[200]=8'he8;
        mem_13[201]=8'hdd;
        mem_13[202]=8'h74;
        mem_13[203]=8'h1f;
        mem_13[204]=8'h4b;
        mem_13[205]=8'hbd;
        mem_13[206]=8'h8b;
        mem_13[207]=8'h8a;
        mem_13[208]=8'h70;
        mem_13[209]=8'h3e;
        mem_13[210]=8'hb5;
        mem_13[211]=8'h66;
        mem_13[212]=8'h48;
        mem_13[213]=8'h3;
        mem_13[214]=8'hf6;
        mem_13[215]=8'he;
        mem_13[216]=8'h61;
        mem_13[217]=8'h35;
        mem_13[218]=8'h57;
        mem_13[219]=8'hb9;
        mem_13[220]=8'h86;
        mem_13[221]=8'hc1;
        mem_13[222]=8'h1d;
        mem_13[223]=8'h9e;
        mem_13[224]=8'he1;
        mem_13[225]=8'hf8;
        mem_13[226]=8'h98;
        mem_13[227]=8'h11;
        mem_13[228]=8'h69;
        mem_13[229]=8'hd9;
        mem_13[230]=8'h8e;
        mem_13[231]=8'h94;
        mem_13[232]=8'h9b;
        mem_13[233]=8'h1e;
        mem_13[234]=8'h87;
        mem_13[235]=8'he9;
        mem_13[236]=8'hce;
        mem_13[237]=8'h55;
        mem_13[238]=8'h28;
        mem_13[239]=8'hdf;
        mem_13[240]=8'h8c;
        mem_13[241]=8'ha1;
        mem_13[242]=8'h89;
        mem_13[243]=8'hd;
        mem_13[244]=8'hbf;
        mem_13[245]=8'he6;
        mem_13[246]=8'h42;
        mem_13[247]=8'h68;
        mem_13[248]=8'h41;
        mem_13[249]=8'h99;
        mem_13[250]=8'h2d;
        mem_13[251]=8'hf;
        mem_13[252]=8'hb0;
        mem_13[253]=8'h54;
        mem_13[254]=8'hbb;
        mem_13[255]=8'h16;
    end

    initial begin
        mem_14[0]=8'h63;
        mem_14[1]=8'h7c;
        mem_14[2]=8'h77;
        mem_14[3]=8'h7b;
        mem_14[4]=8'hf2;
        mem_14[5]=8'h6b;
        mem_14[6]=8'h6f;
        mem_14[7]=8'hc5;
        mem_14[8]=8'h30;
        mem_14[9]=8'h1;
        mem_14[10]=8'h67;
        mem_14[11]=8'h2b;
        mem_14[12]=8'hfe;
        mem_14[13]=8'hd7;
        mem_14[14]=8'hab;
        mem_14[15]=8'h76;
        mem_14[16]=8'hca;
        mem_14[17]=8'h82;
        mem_14[18]=8'hc9;
        mem_14[19]=8'h7d;
        mem_14[20]=8'hfa;
        mem_14[21]=8'h59;
        mem_14[22]=8'h47;
        mem_14[23]=8'hf0;
        mem_14[24]=8'had;
        mem_14[25]=8'hd4;
        mem_14[26]=8'ha2;
        mem_14[27]=8'haf;
        mem_14[28]=8'h9c;
        mem_14[29]=8'ha4;
        mem_14[30]=8'h72;
        mem_14[31]=8'hc0;
        mem_14[32]=8'hb7;
        mem_14[33]=8'hfd;
        mem_14[34]=8'h93;
        mem_14[35]=8'h26;
        mem_14[36]=8'h36;
        mem_14[37]=8'h3f;
        mem_14[38]=8'hf7;
        mem_14[39]=8'hcc;
        mem_14[40]=8'h34;
        mem_14[41]=8'ha5;
        mem_14[42]=8'he5;
        mem_14[43]=8'hf1;
        mem_14[44]=8'h71;
        mem_14[45]=8'hd8;
        mem_14[46]=8'h31;
        mem_14[47]=8'h15;
        mem_14[48]=8'h4;
        mem_14[49]=8'hc7;
        mem_14[50]=8'h23;
        mem_14[51]=8'hc3;
        mem_14[52]=8'h18;
        mem_14[53]=8'h96;
        mem_14[54]=8'h5;
        mem_14[55]=8'h9a;
        mem_14[56]=8'h7;
        mem_14[57]=8'h12;
        mem_14[58]=8'h80;
        mem_14[59]=8'he2;
        mem_14[60]=8'heb;
        mem_14[61]=8'h27;
        mem_14[62]=8'hb2;
        mem_14[63]=8'h75;
        mem_14[64]=8'h9;
        mem_14[65]=8'h83;
        mem_14[66]=8'h2c;
        mem_14[67]=8'h1a;
        mem_14[68]=8'h1b;
        mem_14[69]=8'h6e;
        mem_14[70]=8'h5a;
        mem_14[71]=8'ha0;
        mem_14[72]=8'h52;
        mem_14[73]=8'h3b;
        mem_14[74]=8'hd6;
        mem_14[75]=8'hb3;
        mem_14[76]=8'h29;
        mem_14[77]=8'he3;
        mem_14[78]=8'h2f;
        mem_14[79]=8'h84;
        mem_14[80]=8'h53;
        mem_14[81]=8'hd1;
        mem_14[82]=8'h0;
        mem_14[83]=8'hed;
        mem_14[84]=8'h20;
        mem_14[85]=8'hfc;
        mem_14[86]=8'hb1;
        mem_14[87]=8'h5b;
        mem_14[88]=8'h6a;
        mem_14[89]=8'hcb;
        mem_14[90]=8'hbe;
        mem_14[91]=8'h39;
        mem_14[92]=8'h4a;
        mem_14[93]=8'h4c;
        mem_14[94]=8'h58;
        mem_14[95]=8'hcf;
        mem_14[96]=8'hd0;
        mem_14[97]=8'hef;
        mem_14[98]=8'haa;
        mem_14[99]=8'hfb;
        mem_14[100]=8'h43;
        mem_14[101]=8'h4d;
        mem_14[102]=8'h33;
        mem_14[103]=8'h85;
        mem_14[104]=8'h45;
        mem_14[105]=8'hf9;
        mem_14[106]=8'h2;
        mem_14[107]=8'h7f;
        mem_14[108]=8'h50;
        mem_14[109]=8'h3c;
        mem_14[110]=8'h9f;
        mem_14[111]=8'ha8;
        mem_14[112]=8'h51;
        mem_14[113]=8'ha3;
        mem_14[114]=8'h40;
        mem_14[115]=8'h8f;
        mem_14[116]=8'h92;
        mem_14[117]=8'h9d;
        mem_14[118]=8'h38;
        mem_14[119]=8'hf5;
        mem_14[120]=8'hbc;
        mem_14[121]=8'hb6;
        mem_14[122]=8'hda;
        mem_14[123]=8'h21;
        mem_14[124]=8'h10;
        mem_14[125]=8'hff;
        mem_14[126]=8'hf3;
        mem_14[127]=8'hd2;
        mem_14[128]=8'hcd;
        mem_14[129]=8'hc;
        mem_14[130]=8'h13;
        mem_14[131]=8'hec;
        mem_14[132]=8'h5f;
        mem_14[133]=8'h97;
        mem_14[134]=8'h44;
        mem_14[135]=8'h17;
        mem_14[136]=8'hc4;
        mem_14[137]=8'ha7;
        mem_14[138]=8'h7e;
        mem_14[139]=8'h3d;
        mem_14[140]=8'h64;
        mem_14[141]=8'h5d;
        mem_14[142]=8'h19;
        mem_14[143]=8'h73;
        mem_14[144]=8'h60;
        mem_14[145]=8'h81;
        mem_14[146]=8'h4f;
        mem_14[147]=8'hdc;
        mem_14[148]=8'h22;
        mem_14[149]=8'h2a;
        mem_14[150]=8'h90;
        mem_14[151]=8'h88;
        mem_14[152]=8'h46;
        mem_14[153]=8'hee;
        mem_14[154]=8'hb8;
        mem_14[155]=8'h14;
        mem_14[156]=8'hde;
        mem_14[157]=8'h5e;
        mem_14[158]=8'hb;
        mem_14[159]=8'hdb;
        mem_14[160]=8'he0;
        mem_14[161]=8'h32;
        mem_14[162]=8'h3a;
        mem_14[163]=8'ha;
        mem_14[164]=8'h49;
        mem_14[165]=8'h6;
        mem_14[166]=8'h24;
        mem_14[167]=8'h5c;
        mem_14[168]=8'hc2;
        mem_14[169]=8'hd3;
        mem_14[170]=8'hac;
        mem_14[171]=8'h62;
        mem_14[172]=8'h91;
        mem_14[173]=8'h95;
        mem_14[174]=8'he4;
        mem_14[175]=8'h79;
        mem_14[176]=8'he7;
        mem_14[177]=8'hc8;
        mem_14[178]=8'h37;
        mem_14[179]=8'h6d;
        mem_14[180]=8'h8d;
        mem_14[181]=8'hd5;
        mem_14[182]=8'h4e;
        mem_14[183]=8'ha9;
        mem_14[184]=8'h6c;
        mem_14[185]=8'h56;
        mem_14[186]=8'hf4;
        mem_14[187]=8'hea;
        mem_14[188]=8'h65;
        mem_14[189]=8'h7a;
        mem_14[190]=8'hae;
        mem_14[191]=8'h8;
        mem_14[192]=8'hba;
        mem_14[193]=8'h78;
        mem_14[194]=8'h25;
        mem_14[195]=8'h2e;
        mem_14[196]=8'h1c;
        mem_14[197]=8'ha6;
        mem_14[198]=8'hb4;
        mem_14[199]=8'hc6;
        mem_14[200]=8'he8;
        mem_14[201]=8'hdd;
        mem_14[202]=8'h74;
        mem_14[203]=8'h1f;
        mem_14[204]=8'h4b;
        mem_14[205]=8'hbd;
        mem_14[206]=8'h8b;
        mem_14[207]=8'h8a;
        mem_14[208]=8'h70;
        mem_14[209]=8'h3e;
        mem_14[210]=8'hb5;
        mem_14[211]=8'h66;
        mem_14[212]=8'h48;
        mem_14[213]=8'h3;
        mem_14[214]=8'hf6;
        mem_14[215]=8'he;
        mem_14[216]=8'h61;
        mem_14[217]=8'h35;
        mem_14[218]=8'h57;
        mem_14[219]=8'hb9;
        mem_14[220]=8'h86;
        mem_14[221]=8'hc1;
        mem_14[222]=8'h1d;
        mem_14[223]=8'h9e;
        mem_14[224]=8'he1;
        mem_14[225]=8'hf8;
        mem_14[226]=8'h98;
        mem_14[227]=8'h11;
        mem_14[228]=8'h69;
        mem_14[229]=8'hd9;
        mem_14[230]=8'h8e;
        mem_14[231]=8'h94;
        mem_14[232]=8'h9b;
        mem_14[233]=8'h1e;
        mem_14[234]=8'h87;
        mem_14[235]=8'he9;
        mem_14[236]=8'hce;
        mem_14[237]=8'h55;
        mem_14[238]=8'h28;
        mem_14[239]=8'hdf;
        mem_14[240]=8'h8c;
        mem_14[241]=8'ha1;
        mem_14[242]=8'h89;
        mem_14[243]=8'hd;
        mem_14[244]=8'hbf;
        mem_14[245]=8'he6;
        mem_14[246]=8'h42;
        mem_14[247]=8'h68;
        mem_14[248]=8'h41;
        mem_14[249]=8'h99;
        mem_14[250]=8'h2d;
        mem_14[251]=8'hf;
        mem_14[252]=8'hb0;
        mem_14[253]=8'h54;
        mem_14[254]=8'hbb;
        mem_14[255]=8'h16;
    end

    initial begin
        mem_15[0]=8'h63;
        mem_15[1]=8'h7c;
        mem_15[2]=8'h77;
        mem_15[3]=8'h7b;
        mem_15[4]=8'hf2;
        mem_15[5]=8'h6b;
        mem_15[6]=8'h6f;
        mem_15[7]=8'hc5;
        mem_15[8]=8'h30;
        mem_15[9]=8'h1;
        mem_15[10]=8'h67;
        mem_15[11]=8'h2b;
        mem_15[12]=8'hfe;
        mem_15[13]=8'hd7;
        mem_15[14]=8'hab;
        mem_15[15]=8'h76;
        mem_15[16]=8'hca;
        mem_15[17]=8'h82;
        mem_15[18]=8'hc9;
        mem_15[19]=8'h7d;
        mem_15[20]=8'hfa;
        mem_15[21]=8'h59;
        mem_15[22]=8'h47;
        mem_15[23]=8'hf0;
        mem_15[24]=8'had;
        mem_15[25]=8'hd4;
        mem_15[26]=8'ha2;
        mem_15[27]=8'haf;
        mem_15[28]=8'h9c;
        mem_15[29]=8'ha4;
        mem_15[30]=8'h72;
        mem_15[31]=8'hc0;
        mem_15[32]=8'hb7;
        mem_15[33]=8'hfd;
        mem_15[34]=8'h93;
        mem_15[35]=8'h26;
        mem_15[36]=8'h36;
        mem_15[37]=8'h3f;
        mem_15[38]=8'hf7;
        mem_15[39]=8'hcc;
        mem_15[40]=8'h34;
        mem_15[41]=8'ha5;
        mem_15[42]=8'he5;
        mem_15[43]=8'hf1;
        mem_15[44]=8'h71;
        mem_15[45]=8'hd8;
        mem_15[46]=8'h31;
        mem_15[47]=8'h15;
        mem_15[48]=8'h4;
        mem_15[49]=8'hc7;
        mem_15[50]=8'h23;
        mem_15[51]=8'hc3;
        mem_15[52]=8'h18;
        mem_15[53]=8'h96;
        mem_15[54]=8'h5;
        mem_15[55]=8'h9a;
        mem_15[56]=8'h7;
        mem_15[57]=8'h12;
        mem_15[58]=8'h80;
        mem_15[59]=8'he2;
        mem_15[60]=8'heb;
        mem_15[61]=8'h27;
        mem_15[62]=8'hb2;
        mem_15[63]=8'h75;
        mem_15[64]=8'h9;
        mem_15[65]=8'h83;
        mem_15[66]=8'h2c;
        mem_15[67]=8'h1a;
        mem_15[68]=8'h1b;
        mem_15[69]=8'h6e;
        mem_15[70]=8'h5a;
        mem_15[71]=8'ha0;
        mem_15[72]=8'h52;
        mem_15[73]=8'h3b;
        mem_15[74]=8'hd6;
        mem_15[75]=8'hb3;
        mem_15[76]=8'h29;
        mem_15[77]=8'he3;
        mem_15[78]=8'h2f;
        mem_15[79]=8'h84;
        mem_15[80]=8'h53;
        mem_15[81]=8'hd1;
        mem_15[82]=8'h0;
        mem_15[83]=8'hed;
        mem_15[84]=8'h20;
        mem_15[85]=8'hfc;
        mem_15[86]=8'hb1;
        mem_15[87]=8'h5b;
        mem_15[88]=8'h6a;
        mem_15[89]=8'hcb;
        mem_15[90]=8'hbe;
        mem_15[91]=8'h39;
        mem_15[92]=8'h4a;
        mem_15[93]=8'h4c;
        mem_15[94]=8'h58;
        mem_15[95]=8'hcf;
        mem_15[96]=8'hd0;
        mem_15[97]=8'hef;
        mem_15[98]=8'haa;
        mem_15[99]=8'hfb;
        mem_15[100]=8'h43;
        mem_15[101]=8'h4d;
        mem_15[102]=8'h33;
        mem_15[103]=8'h85;
        mem_15[104]=8'h45;
        mem_15[105]=8'hf9;
        mem_15[106]=8'h2;
        mem_15[107]=8'h7f;
        mem_15[108]=8'h50;
        mem_15[109]=8'h3c;
        mem_15[110]=8'h9f;
        mem_15[111]=8'ha8;
        mem_15[112]=8'h51;
        mem_15[113]=8'ha3;
        mem_15[114]=8'h40;
        mem_15[115]=8'h8f;
        mem_15[116]=8'h92;
        mem_15[117]=8'h9d;
        mem_15[118]=8'h38;
        mem_15[119]=8'hf5;
        mem_15[120]=8'hbc;
        mem_15[121]=8'hb6;
        mem_15[122]=8'hda;
        mem_15[123]=8'h21;
        mem_15[124]=8'h10;
        mem_15[125]=8'hff;
        mem_15[126]=8'hf3;
        mem_15[127]=8'hd2;
        mem_15[128]=8'hcd;
        mem_15[129]=8'hc;
        mem_15[130]=8'h13;
        mem_15[131]=8'hec;
        mem_15[132]=8'h5f;
        mem_15[133]=8'h97;
        mem_15[134]=8'h44;
        mem_15[135]=8'h17;
        mem_15[136]=8'hc4;
        mem_15[137]=8'ha7;
        mem_15[138]=8'h7e;
        mem_15[139]=8'h3d;
        mem_15[140]=8'h64;
        mem_15[141]=8'h5d;
        mem_15[142]=8'h19;
        mem_15[143]=8'h73;
        mem_15[144]=8'h60;
        mem_15[145]=8'h81;
        mem_15[146]=8'h4f;
        mem_15[147]=8'hdc;
        mem_15[148]=8'h22;
        mem_15[149]=8'h2a;
        mem_15[150]=8'h90;
        mem_15[151]=8'h88;
        mem_15[152]=8'h46;
        mem_15[153]=8'hee;
        mem_15[154]=8'hb8;
        mem_15[155]=8'h14;
        mem_15[156]=8'hde;
        mem_15[157]=8'h5e;
        mem_15[158]=8'hb;
        mem_15[159]=8'hdb;
        mem_15[160]=8'he0;
        mem_15[161]=8'h32;
        mem_15[162]=8'h3a;
        mem_15[163]=8'ha;
        mem_15[164]=8'h49;
        mem_15[165]=8'h6;
        mem_15[166]=8'h24;
        mem_15[167]=8'h5c;
        mem_15[168]=8'hc2;
        mem_15[169]=8'hd3;
        mem_15[170]=8'hac;
        mem_15[171]=8'h62;
        mem_15[172]=8'h91;
        mem_15[173]=8'h95;
        mem_15[174]=8'he4;
        mem_15[175]=8'h79;
        mem_15[176]=8'he7;
        mem_15[177]=8'hc8;
        mem_15[178]=8'h37;
        mem_15[179]=8'h6d;
        mem_15[180]=8'h8d;
        mem_15[181]=8'hd5;
        mem_15[182]=8'h4e;
        mem_15[183]=8'ha9;
        mem_15[184]=8'h6c;
        mem_15[185]=8'h56;
        mem_15[186]=8'hf4;
        mem_15[187]=8'hea;
        mem_15[188]=8'h65;
        mem_15[189]=8'h7a;
        mem_15[190]=8'hae;
        mem_15[191]=8'h8;
        mem_15[192]=8'hba;
        mem_15[193]=8'h78;
        mem_15[194]=8'h25;
        mem_15[195]=8'h2e;
        mem_15[196]=8'h1c;
        mem_15[197]=8'ha6;
        mem_15[198]=8'hb4;
        mem_15[199]=8'hc6;
        mem_15[200]=8'he8;
        mem_15[201]=8'hdd;
        mem_15[202]=8'h74;
        mem_15[203]=8'h1f;
        mem_15[204]=8'h4b;
        mem_15[205]=8'hbd;
        mem_15[206]=8'h8b;
        mem_15[207]=8'h8a;
        mem_15[208]=8'h70;
        mem_15[209]=8'h3e;
        mem_15[210]=8'hb5;
        mem_15[211]=8'h66;
        mem_15[212]=8'h48;
        mem_15[213]=8'h3;
        mem_15[214]=8'hf6;
        mem_15[215]=8'he;
        mem_15[216]=8'h61;
        mem_15[217]=8'h35;
        mem_15[218]=8'h57;
        mem_15[219]=8'hb9;
        mem_15[220]=8'h86;
        mem_15[221]=8'hc1;
        mem_15[222]=8'h1d;
        mem_15[223]=8'h9e;
        mem_15[224]=8'he1;
        mem_15[225]=8'hf8;
        mem_15[226]=8'h98;
        mem_15[227]=8'h11;
        mem_15[228]=8'h69;
        mem_15[229]=8'hd9;
        mem_15[230]=8'h8e;
        mem_15[231]=8'h94;
        mem_15[232]=8'h9b;
        mem_15[233]=8'h1e;
        mem_15[234]=8'h87;
        mem_15[235]=8'he9;
        mem_15[236]=8'hce;
        mem_15[237]=8'h55;
        mem_15[238]=8'h28;
        mem_15[239]=8'hdf;
        mem_15[240]=8'h8c;
        mem_15[241]=8'ha1;
        mem_15[242]=8'h89;
        mem_15[243]=8'hd;
        mem_15[244]=8'hbf;
        mem_15[245]=8'he6;
        mem_15[246]=8'h42;
        mem_15[247]=8'h68;
        mem_15[248]=8'h41;
        mem_15[249]=8'h99;
        mem_15[250]=8'h2d;
        mem_15[251]=8'hf;
        mem_15[252]=8'hb0;
        mem_15[253]=8'h54;
        mem_15[254]=8'hbb;
        mem_15[255]=8'h16;
    end

    initial begin
        mem_16[0]=8'h63;
        mem_16[1]=8'h7c;
        mem_16[2]=8'h77;
        mem_16[3]=8'h7b;
        mem_16[4]=8'hf2;
        mem_16[5]=8'h6b;
        mem_16[6]=8'h6f;
        mem_16[7]=8'hc5;
        mem_16[8]=8'h30;
        mem_16[9]=8'h1;
        mem_16[10]=8'h67;
        mem_16[11]=8'h2b;
        mem_16[12]=8'hfe;
        mem_16[13]=8'hd7;
        mem_16[14]=8'hab;
        mem_16[15]=8'h76;
        mem_16[16]=8'hca;
        mem_16[17]=8'h82;
        mem_16[18]=8'hc9;
        mem_16[19]=8'h7d;
        mem_16[20]=8'hfa;
        mem_16[21]=8'h59;
        mem_16[22]=8'h47;
        mem_16[23]=8'hf0;
        mem_16[24]=8'had;
        mem_16[25]=8'hd4;
        mem_16[26]=8'ha2;
        mem_16[27]=8'haf;
        mem_16[28]=8'h9c;
        mem_16[29]=8'ha4;
        mem_16[30]=8'h72;
        mem_16[31]=8'hc0;
        mem_16[32]=8'hb7;
        mem_16[33]=8'hfd;
        mem_16[34]=8'h93;
        mem_16[35]=8'h26;
        mem_16[36]=8'h36;
        mem_16[37]=8'h3f;
        mem_16[38]=8'hf7;
        mem_16[39]=8'hcc;
        mem_16[40]=8'h34;
        mem_16[41]=8'ha5;
        mem_16[42]=8'he5;
        mem_16[43]=8'hf1;
        mem_16[44]=8'h71;
        mem_16[45]=8'hd8;
        mem_16[46]=8'h31;
        mem_16[47]=8'h15;
        mem_16[48]=8'h4;
        mem_16[49]=8'hc7;
        mem_16[50]=8'h23;
        mem_16[51]=8'hc3;
        mem_16[52]=8'h18;
        mem_16[53]=8'h96;
        mem_16[54]=8'h5;
        mem_16[55]=8'h9a;
        mem_16[56]=8'h7;
        mem_16[57]=8'h12;
        mem_16[58]=8'h80;
        mem_16[59]=8'he2;
        mem_16[60]=8'heb;
        mem_16[61]=8'h27;
        mem_16[62]=8'hb2;
        mem_16[63]=8'h75;
        mem_16[64]=8'h9;
        mem_16[65]=8'h83;
        mem_16[66]=8'h2c;
        mem_16[67]=8'h1a;
        mem_16[68]=8'h1b;
        mem_16[69]=8'h6e;
        mem_16[70]=8'h5a;
        mem_16[71]=8'ha0;
        mem_16[72]=8'h52;
        mem_16[73]=8'h3b;
        mem_16[74]=8'hd6;
        mem_16[75]=8'hb3;
        mem_16[76]=8'h29;
        mem_16[77]=8'he3;
        mem_16[78]=8'h2f;
        mem_16[79]=8'h84;
        mem_16[80]=8'h53;
        mem_16[81]=8'hd1;
        mem_16[82]=8'h0;
        mem_16[83]=8'hed;
        mem_16[84]=8'h20;
        mem_16[85]=8'hfc;
        mem_16[86]=8'hb1;
        mem_16[87]=8'h5b;
        mem_16[88]=8'h6a;
        mem_16[89]=8'hcb;
        mem_16[90]=8'hbe;
        mem_16[91]=8'h39;
        mem_16[92]=8'h4a;
        mem_16[93]=8'h4c;
        mem_16[94]=8'h58;
        mem_16[95]=8'hcf;
        mem_16[96]=8'hd0;
        mem_16[97]=8'hef;
        mem_16[98]=8'haa;
        mem_16[99]=8'hfb;
        mem_16[100]=8'h43;
        mem_16[101]=8'h4d;
        mem_16[102]=8'h33;
        mem_16[103]=8'h85;
        mem_16[104]=8'h45;
        mem_16[105]=8'hf9;
        mem_16[106]=8'h2;
        mem_16[107]=8'h7f;
        mem_16[108]=8'h50;
        mem_16[109]=8'h3c;
        mem_16[110]=8'h9f;
        mem_16[111]=8'ha8;
        mem_16[112]=8'h51;
        mem_16[113]=8'ha3;
        mem_16[114]=8'h40;
        mem_16[115]=8'h8f;
        mem_16[116]=8'h92;
        mem_16[117]=8'h9d;
        mem_16[118]=8'h38;
        mem_16[119]=8'hf5;
        mem_16[120]=8'hbc;
        mem_16[121]=8'hb6;
        mem_16[122]=8'hda;
        mem_16[123]=8'h21;
        mem_16[124]=8'h10;
        mem_16[125]=8'hff;
        mem_16[126]=8'hf3;
        mem_16[127]=8'hd2;
        mem_16[128]=8'hcd;
        mem_16[129]=8'hc;
        mem_16[130]=8'h13;
        mem_16[131]=8'hec;
        mem_16[132]=8'h5f;
        mem_16[133]=8'h97;
        mem_16[134]=8'h44;
        mem_16[135]=8'h17;
        mem_16[136]=8'hc4;
        mem_16[137]=8'ha7;
        mem_16[138]=8'h7e;
        mem_16[139]=8'h3d;
        mem_16[140]=8'h64;
        mem_16[141]=8'h5d;
        mem_16[142]=8'h19;
        mem_16[143]=8'h73;
        mem_16[144]=8'h60;
        mem_16[145]=8'h81;
        mem_16[146]=8'h4f;
        mem_16[147]=8'hdc;
        mem_16[148]=8'h22;
        mem_16[149]=8'h2a;
        mem_16[150]=8'h90;
        mem_16[151]=8'h88;
        mem_16[152]=8'h46;
        mem_16[153]=8'hee;
        mem_16[154]=8'hb8;
        mem_16[155]=8'h14;
        mem_16[156]=8'hde;
        mem_16[157]=8'h5e;
        mem_16[158]=8'hb;
        mem_16[159]=8'hdb;
        mem_16[160]=8'he0;
        mem_16[161]=8'h32;
        mem_16[162]=8'h3a;
        mem_16[163]=8'ha;
        mem_16[164]=8'h49;
        mem_16[165]=8'h6;
        mem_16[166]=8'h24;
        mem_16[167]=8'h5c;
        mem_16[168]=8'hc2;
        mem_16[169]=8'hd3;
        mem_16[170]=8'hac;
        mem_16[171]=8'h62;
        mem_16[172]=8'h91;
        mem_16[173]=8'h95;
        mem_16[174]=8'he4;
        mem_16[175]=8'h79;
        mem_16[176]=8'he7;
        mem_16[177]=8'hc8;
        mem_16[178]=8'h37;
        mem_16[179]=8'h6d;
        mem_16[180]=8'h8d;
        mem_16[181]=8'hd5;
        mem_16[182]=8'h4e;
        mem_16[183]=8'ha9;
        mem_16[184]=8'h6c;
        mem_16[185]=8'h56;
        mem_16[186]=8'hf4;
        mem_16[187]=8'hea;
        mem_16[188]=8'h65;
        mem_16[189]=8'h7a;
        mem_16[190]=8'hae;
        mem_16[191]=8'h8;
        mem_16[192]=8'hba;
        mem_16[193]=8'h78;
        mem_16[194]=8'h25;
        mem_16[195]=8'h2e;
        mem_16[196]=8'h1c;
        mem_16[197]=8'ha6;
        mem_16[198]=8'hb4;
        mem_16[199]=8'hc6;
        mem_16[200]=8'he8;
        mem_16[201]=8'hdd;
        mem_16[202]=8'h74;
        mem_16[203]=8'h1f;
        mem_16[204]=8'h4b;
        mem_16[205]=8'hbd;
        mem_16[206]=8'h8b;
        mem_16[207]=8'h8a;
        mem_16[208]=8'h70;
        mem_16[209]=8'h3e;
        mem_16[210]=8'hb5;
        mem_16[211]=8'h66;
        mem_16[212]=8'h48;
        mem_16[213]=8'h3;
        mem_16[214]=8'hf6;
        mem_16[215]=8'he;
        mem_16[216]=8'h61;
        mem_16[217]=8'h35;
        mem_16[218]=8'h57;
        mem_16[219]=8'hb9;
        mem_16[220]=8'h86;
        mem_16[221]=8'hc1;
        mem_16[222]=8'h1d;
        mem_16[223]=8'h9e;
        mem_16[224]=8'he1;
        mem_16[225]=8'hf8;
        mem_16[226]=8'h98;
        mem_16[227]=8'h11;
        mem_16[228]=8'h69;
        mem_16[229]=8'hd9;
        mem_16[230]=8'h8e;
        mem_16[231]=8'h94;
        mem_16[232]=8'h9b;
        mem_16[233]=8'h1e;
        mem_16[234]=8'h87;
        mem_16[235]=8'he9;
        mem_16[236]=8'hce;
        mem_16[237]=8'h55;
        mem_16[238]=8'h28;
        mem_16[239]=8'hdf;
        mem_16[240]=8'h8c;
        mem_16[241]=8'ha1;
        mem_16[242]=8'h89;
        mem_16[243]=8'hd;
        mem_16[244]=8'hbf;
        mem_16[245]=8'he6;
        mem_16[246]=8'h42;
        mem_16[247]=8'h68;
        mem_16[248]=8'h41;
        mem_16[249]=8'h99;
        mem_16[250]=8'h2d;
        mem_16[251]=8'hf;
        mem_16[252]=8'hb0;
        mem_16[253]=8'h54;
        mem_16[254]=8'hbb;
        mem_16[255]=8'h16;
    end

    initial begin
        mem_17[0]=8'h63;
        mem_17[1]=8'h7c;
        mem_17[2]=8'h77;
        mem_17[3]=8'h7b;
        mem_17[4]=8'hf2;
        mem_17[5]=8'h6b;
        mem_17[6]=8'h6f;
        mem_17[7]=8'hc5;
        mem_17[8]=8'h30;
        mem_17[9]=8'h1;
        mem_17[10]=8'h67;
        mem_17[11]=8'h2b;
        mem_17[12]=8'hfe;
        mem_17[13]=8'hd7;
        mem_17[14]=8'hab;
        mem_17[15]=8'h76;
        mem_17[16]=8'hca;
        mem_17[17]=8'h82;
        mem_17[18]=8'hc9;
        mem_17[19]=8'h7d;
        mem_17[20]=8'hfa;
        mem_17[21]=8'h59;
        mem_17[22]=8'h47;
        mem_17[23]=8'hf0;
        mem_17[24]=8'had;
        mem_17[25]=8'hd4;
        mem_17[26]=8'ha2;
        mem_17[27]=8'haf;
        mem_17[28]=8'h9c;
        mem_17[29]=8'ha4;
        mem_17[30]=8'h72;
        mem_17[31]=8'hc0;
        mem_17[32]=8'hb7;
        mem_17[33]=8'hfd;
        mem_17[34]=8'h93;
        mem_17[35]=8'h26;
        mem_17[36]=8'h36;
        mem_17[37]=8'h3f;
        mem_17[38]=8'hf7;
        mem_17[39]=8'hcc;
        mem_17[40]=8'h34;
        mem_17[41]=8'ha5;
        mem_17[42]=8'he5;
        mem_17[43]=8'hf1;
        mem_17[44]=8'h71;
        mem_17[45]=8'hd8;
        mem_17[46]=8'h31;
        mem_17[47]=8'h15;
        mem_17[48]=8'h4;
        mem_17[49]=8'hc7;
        mem_17[50]=8'h23;
        mem_17[51]=8'hc3;
        mem_17[52]=8'h18;
        mem_17[53]=8'h96;
        mem_17[54]=8'h5;
        mem_17[55]=8'h9a;
        mem_17[56]=8'h7;
        mem_17[57]=8'h12;
        mem_17[58]=8'h80;
        mem_17[59]=8'he2;
        mem_17[60]=8'heb;
        mem_17[61]=8'h27;
        mem_17[62]=8'hb2;
        mem_17[63]=8'h75;
        mem_17[64]=8'h9;
        mem_17[65]=8'h83;
        mem_17[66]=8'h2c;
        mem_17[67]=8'h1a;
        mem_17[68]=8'h1b;
        mem_17[69]=8'h6e;
        mem_17[70]=8'h5a;
        mem_17[71]=8'ha0;
        mem_17[72]=8'h52;
        mem_17[73]=8'h3b;
        mem_17[74]=8'hd6;
        mem_17[75]=8'hb3;
        mem_17[76]=8'h29;
        mem_17[77]=8'he3;
        mem_17[78]=8'h2f;
        mem_17[79]=8'h84;
        mem_17[80]=8'h53;
        mem_17[81]=8'hd1;
        mem_17[82]=8'h0;
        mem_17[83]=8'hed;
        mem_17[84]=8'h20;
        mem_17[85]=8'hfc;
        mem_17[86]=8'hb1;
        mem_17[87]=8'h5b;
        mem_17[88]=8'h6a;
        mem_17[89]=8'hcb;
        mem_17[90]=8'hbe;
        mem_17[91]=8'h39;
        mem_17[92]=8'h4a;
        mem_17[93]=8'h4c;
        mem_17[94]=8'h58;
        mem_17[95]=8'hcf;
        mem_17[96]=8'hd0;
        mem_17[97]=8'hef;
        mem_17[98]=8'haa;
        mem_17[99]=8'hfb;
        mem_17[100]=8'h43;
        mem_17[101]=8'h4d;
        mem_17[102]=8'h33;
        mem_17[103]=8'h85;
        mem_17[104]=8'h45;
        mem_17[105]=8'hf9;
        mem_17[106]=8'h2;
        mem_17[107]=8'h7f;
        mem_17[108]=8'h50;
        mem_17[109]=8'h3c;
        mem_17[110]=8'h9f;
        mem_17[111]=8'ha8;
        mem_17[112]=8'h51;
        mem_17[113]=8'ha3;
        mem_17[114]=8'h40;
        mem_17[115]=8'h8f;
        mem_17[116]=8'h92;
        mem_17[117]=8'h9d;
        mem_17[118]=8'h38;
        mem_17[119]=8'hf5;
        mem_17[120]=8'hbc;
        mem_17[121]=8'hb6;
        mem_17[122]=8'hda;
        mem_17[123]=8'h21;
        mem_17[124]=8'h10;
        mem_17[125]=8'hff;
        mem_17[126]=8'hf3;
        mem_17[127]=8'hd2;
        mem_17[128]=8'hcd;
        mem_17[129]=8'hc;
        mem_17[130]=8'h13;
        mem_17[131]=8'hec;
        mem_17[132]=8'h5f;
        mem_17[133]=8'h97;
        mem_17[134]=8'h44;
        mem_17[135]=8'h17;
        mem_17[136]=8'hc4;
        mem_17[137]=8'ha7;
        mem_17[138]=8'h7e;
        mem_17[139]=8'h3d;
        mem_17[140]=8'h64;
        mem_17[141]=8'h5d;
        mem_17[142]=8'h19;
        mem_17[143]=8'h73;
        mem_17[144]=8'h60;
        mem_17[145]=8'h81;
        mem_17[146]=8'h4f;
        mem_17[147]=8'hdc;
        mem_17[148]=8'h22;
        mem_17[149]=8'h2a;
        mem_17[150]=8'h90;
        mem_17[151]=8'h88;
        mem_17[152]=8'h46;
        mem_17[153]=8'hee;
        mem_17[154]=8'hb8;
        mem_17[155]=8'h14;
        mem_17[156]=8'hde;
        mem_17[157]=8'h5e;
        mem_17[158]=8'hb;
        mem_17[159]=8'hdb;
        mem_17[160]=8'he0;
        mem_17[161]=8'h32;
        mem_17[162]=8'h3a;
        mem_17[163]=8'ha;
        mem_17[164]=8'h49;
        mem_17[165]=8'h6;
        mem_17[166]=8'h24;
        mem_17[167]=8'h5c;
        mem_17[168]=8'hc2;
        mem_17[169]=8'hd3;
        mem_17[170]=8'hac;
        mem_17[171]=8'h62;
        mem_17[172]=8'h91;
        mem_17[173]=8'h95;
        mem_17[174]=8'he4;
        mem_17[175]=8'h79;
        mem_17[176]=8'he7;
        mem_17[177]=8'hc8;
        mem_17[178]=8'h37;
        mem_17[179]=8'h6d;
        mem_17[180]=8'h8d;
        mem_17[181]=8'hd5;
        mem_17[182]=8'h4e;
        mem_17[183]=8'ha9;
        mem_17[184]=8'h6c;
        mem_17[185]=8'h56;
        mem_17[186]=8'hf4;
        mem_17[187]=8'hea;
        mem_17[188]=8'h65;
        mem_17[189]=8'h7a;
        mem_17[190]=8'hae;
        mem_17[191]=8'h8;
        mem_17[192]=8'hba;
        mem_17[193]=8'h78;
        mem_17[194]=8'h25;
        mem_17[195]=8'h2e;
        mem_17[196]=8'h1c;
        mem_17[197]=8'ha6;
        mem_17[198]=8'hb4;
        mem_17[199]=8'hc6;
        mem_17[200]=8'he8;
        mem_17[201]=8'hdd;
        mem_17[202]=8'h74;
        mem_17[203]=8'h1f;
        mem_17[204]=8'h4b;
        mem_17[205]=8'hbd;
        mem_17[206]=8'h8b;
        mem_17[207]=8'h8a;
        mem_17[208]=8'h70;
        mem_17[209]=8'h3e;
        mem_17[210]=8'hb5;
        mem_17[211]=8'h66;
        mem_17[212]=8'h48;
        mem_17[213]=8'h3;
        mem_17[214]=8'hf6;
        mem_17[215]=8'he;
        mem_17[216]=8'h61;
        mem_17[217]=8'h35;
        mem_17[218]=8'h57;
        mem_17[219]=8'hb9;
        mem_17[220]=8'h86;
        mem_17[221]=8'hc1;
        mem_17[222]=8'h1d;
        mem_17[223]=8'h9e;
        mem_17[224]=8'he1;
        mem_17[225]=8'hf8;
        mem_17[226]=8'h98;
        mem_17[227]=8'h11;
        mem_17[228]=8'h69;
        mem_17[229]=8'hd9;
        mem_17[230]=8'h8e;
        mem_17[231]=8'h94;
        mem_17[232]=8'h9b;
        mem_17[233]=8'h1e;
        mem_17[234]=8'h87;
        mem_17[235]=8'he9;
        mem_17[236]=8'hce;
        mem_17[237]=8'h55;
        mem_17[238]=8'h28;
        mem_17[239]=8'hdf;
        mem_17[240]=8'h8c;
        mem_17[241]=8'ha1;
        mem_17[242]=8'h89;
        mem_17[243]=8'hd;
        mem_17[244]=8'hbf;
        mem_17[245]=8'he6;
        mem_17[246]=8'h42;
        mem_17[247]=8'h68;
        mem_17[248]=8'h41;
        mem_17[249]=8'h99;
        mem_17[250]=8'h2d;
        mem_17[251]=8'hf;
        mem_17[252]=8'hb0;
        mem_17[253]=8'h54;
        mem_17[254]=8'hbb;
        mem_17[255]=8'h16;
    end

    initial begin
        mem_18[0]=8'h63;
        mem_18[1]=8'h7c;
        mem_18[2]=8'h77;
        mem_18[3]=8'h7b;
        mem_18[4]=8'hf2;
        mem_18[5]=8'h6b;
        mem_18[6]=8'h6f;
        mem_18[7]=8'hc5;
        mem_18[8]=8'h30;
        mem_18[9]=8'h1;
        mem_18[10]=8'h67;
        mem_18[11]=8'h2b;
        mem_18[12]=8'hfe;
        mem_18[13]=8'hd7;
        mem_18[14]=8'hab;
        mem_18[15]=8'h76;
        mem_18[16]=8'hca;
        mem_18[17]=8'h82;
        mem_18[18]=8'hc9;
        mem_18[19]=8'h7d;
        mem_18[20]=8'hfa;
        mem_18[21]=8'h59;
        mem_18[22]=8'h47;
        mem_18[23]=8'hf0;
        mem_18[24]=8'had;
        mem_18[25]=8'hd4;
        mem_18[26]=8'ha2;
        mem_18[27]=8'haf;
        mem_18[28]=8'h9c;
        mem_18[29]=8'ha4;
        mem_18[30]=8'h72;
        mem_18[31]=8'hc0;
        mem_18[32]=8'hb7;
        mem_18[33]=8'hfd;
        mem_18[34]=8'h93;
        mem_18[35]=8'h26;
        mem_18[36]=8'h36;
        mem_18[37]=8'h3f;
        mem_18[38]=8'hf7;
        mem_18[39]=8'hcc;
        mem_18[40]=8'h34;
        mem_18[41]=8'ha5;
        mem_18[42]=8'he5;
        mem_18[43]=8'hf1;
        mem_18[44]=8'h71;
        mem_18[45]=8'hd8;
        mem_18[46]=8'h31;
        mem_18[47]=8'h15;
        mem_18[48]=8'h4;
        mem_18[49]=8'hc7;
        mem_18[50]=8'h23;
        mem_18[51]=8'hc3;
        mem_18[52]=8'h18;
        mem_18[53]=8'h96;
        mem_18[54]=8'h5;
        mem_18[55]=8'h9a;
        mem_18[56]=8'h7;
        mem_18[57]=8'h12;
        mem_18[58]=8'h80;
        mem_18[59]=8'he2;
        mem_18[60]=8'heb;
        mem_18[61]=8'h27;
        mem_18[62]=8'hb2;
        mem_18[63]=8'h75;
        mem_18[64]=8'h9;
        mem_18[65]=8'h83;
        mem_18[66]=8'h2c;
        mem_18[67]=8'h1a;
        mem_18[68]=8'h1b;
        mem_18[69]=8'h6e;
        mem_18[70]=8'h5a;
        mem_18[71]=8'ha0;
        mem_18[72]=8'h52;
        mem_18[73]=8'h3b;
        mem_18[74]=8'hd6;
        mem_18[75]=8'hb3;
        mem_18[76]=8'h29;
        mem_18[77]=8'he3;
        mem_18[78]=8'h2f;
        mem_18[79]=8'h84;
        mem_18[80]=8'h53;
        mem_18[81]=8'hd1;
        mem_18[82]=8'h0;
        mem_18[83]=8'hed;
        mem_18[84]=8'h20;
        mem_18[85]=8'hfc;
        mem_18[86]=8'hb1;
        mem_18[87]=8'h5b;
        mem_18[88]=8'h6a;
        mem_18[89]=8'hcb;
        mem_18[90]=8'hbe;
        mem_18[91]=8'h39;
        mem_18[92]=8'h4a;
        mem_18[93]=8'h4c;
        mem_18[94]=8'h58;
        mem_18[95]=8'hcf;
        mem_18[96]=8'hd0;
        mem_18[97]=8'hef;
        mem_18[98]=8'haa;
        mem_18[99]=8'hfb;
        mem_18[100]=8'h43;
        mem_18[101]=8'h4d;
        mem_18[102]=8'h33;
        mem_18[103]=8'h85;
        mem_18[104]=8'h45;
        mem_18[105]=8'hf9;
        mem_18[106]=8'h2;
        mem_18[107]=8'h7f;
        mem_18[108]=8'h50;
        mem_18[109]=8'h3c;
        mem_18[110]=8'h9f;
        mem_18[111]=8'ha8;
        mem_18[112]=8'h51;
        mem_18[113]=8'ha3;
        mem_18[114]=8'h40;
        mem_18[115]=8'h8f;
        mem_18[116]=8'h92;
        mem_18[117]=8'h9d;
        mem_18[118]=8'h38;
        mem_18[119]=8'hf5;
        mem_18[120]=8'hbc;
        mem_18[121]=8'hb6;
        mem_18[122]=8'hda;
        mem_18[123]=8'h21;
        mem_18[124]=8'h10;
        mem_18[125]=8'hff;
        mem_18[126]=8'hf3;
        mem_18[127]=8'hd2;
        mem_18[128]=8'hcd;
        mem_18[129]=8'hc;
        mem_18[130]=8'h13;
        mem_18[131]=8'hec;
        mem_18[132]=8'h5f;
        mem_18[133]=8'h97;
        mem_18[134]=8'h44;
        mem_18[135]=8'h17;
        mem_18[136]=8'hc4;
        mem_18[137]=8'ha7;
        mem_18[138]=8'h7e;
        mem_18[139]=8'h3d;
        mem_18[140]=8'h64;
        mem_18[141]=8'h5d;
        mem_18[142]=8'h19;
        mem_18[143]=8'h73;
        mem_18[144]=8'h60;
        mem_18[145]=8'h81;
        mem_18[146]=8'h4f;
        mem_18[147]=8'hdc;
        mem_18[148]=8'h22;
        mem_18[149]=8'h2a;
        mem_18[150]=8'h90;
        mem_18[151]=8'h88;
        mem_18[152]=8'h46;
        mem_18[153]=8'hee;
        mem_18[154]=8'hb8;
        mem_18[155]=8'h14;
        mem_18[156]=8'hde;
        mem_18[157]=8'h5e;
        mem_18[158]=8'hb;
        mem_18[159]=8'hdb;
        mem_18[160]=8'he0;
        mem_18[161]=8'h32;
        mem_18[162]=8'h3a;
        mem_18[163]=8'ha;
        mem_18[164]=8'h49;
        mem_18[165]=8'h6;
        mem_18[166]=8'h24;
        mem_18[167]=8'h5c;
        mem_18[168]=8'hc2;
        mem_18[169]=8'hd3;
        mem_18[170]=8'hac;
        mem_18[171]=8'h62;
        mem_18[172]=8'h91;
        mem_18[173]=8'h95;
        mem_18[174]=8'he4;
        mem_18[175]=8'h79;
        mem_18[176]=8'he7;
        mem_18[177]=8'hc8;
        mem_18[178]=8'h37;
        mem_18[179]=8'h6d;
        mem_18[180]=8'h8d;
        mem_18[181]=8'hd5;
        mem_18[182]=8'h4e;
        mem_18[183]=8'ha9;
        mem_18[184]=8'h6c;
        mem_18[185]=8'h56;
        mem_18[186]=8'hf4;
        mem_18[187]=8'hea;
        mem_18[188]=8'h65;
        mem_18[189]=8'h7a;
        mem_18[190]=8'hae;
        mem_18[191]=8'h8;
        mem_18[192]=8'hba;
        mem_18[193]=8'h78;
        mem_18[194]=8'h25;
        mem_18[195]=8'h2e;
        mem_18[196]=8'h1c;
        mem_18[197]=8'ha6;
        mem_18[198]=8'hb4;
        mem_18[199]=8'hc6;
        mem_18[200]=8'he8;
        mem_18[201]=8'hdd;
        mem_18[202]=8'h74;
        mem_18[203]=8'h1f;
        mem_18[204]=8'h4b;
        mem_18[205]=8'hbd;
        mem_18[206]=8'h8b;
        mem_18[207]=8'h8a;
        mem_18[208]=8'h70;
        mem_18[209]=8'h3e;
        mem_18[210]=8'hb5;
        mem_18[211]=8'h66;
        mem_18[212]=8'h48;
        mem_18[213]=8'h3;
        mem_18[214]=8'hf6;
        mem_18[215]=8'he;
        mem_18[216]=8'h61;
        mem_18[217]=8'h35;
        mem_18[218]=8'h57;
        mem_18[219]=8'hb9;
        mem_18[220]=8'h86;
        mem_18[221]=8'hc1;
        mem_18[222]=8'h1d;
        mem_18[223]=8'h9e;
        mem_18[224]=8'he1;
        mem_18[225]=8'hf8;
        mem_18[226]=8'h98;
        mem_18[227]=8'h11;
        mem_18[228]=8'h69;
        mem_18[229]=8'hd9;
        mem_18[230]=8'h8e;
        mem_18[231]=8'h94;
        mem_18[232]=8'h9b;
        mem_18[233]=8'h1e;
        mem_18[234]=8'h87;
        mem_18[235]=8'he9;
        mem_18[236]=8'hce;
        mem_18[237]=8'h55;
        mem_18[238]=8'h28;
        mem_18[239]=8'hdf;
        mem_18[240]=8'h8c;
        mem_18[241]=8'ha1;
        mem_18[242]=8'h89;
        mem_18[243]=8'hd;
        mem_18[244]=8'hbf;
        mem_18[245]=8'he6;
        mem_18[246]=8'h42;
        mem_18[247]=8'h68;
        mem_18[248]=8'h41;
        mem_18[249]=8'h99;
        mem_18[250]=8'h2d;
        mem_18[251]=8'hf;
        mem_18[252]=8'hb0;
        mem_18[253]=8'h54;
        mem_18[254]=8'hbb;
        mem_18[255]=8'h16;
    end

    initial begin
        mem_19[0]=8'h63;
        mem_19[1]=8'h7c;
        mem_19[2]=8'h77;
        mem_19[3]=8'h7b;
        mem_19[4]=8'hf2;
        mem_19[5]=8'h6b;
        mem_19[6]=8'h6f;
        mem_19[7]=8'hc5;
        mem_19[8]=8'h30;
        mem_19[9]=8'h1;
        mem_19[10]=8'h67;
        mem_19[11]=8'h2b;
        mem_19[12]=8'hfe;
        mem_19[13]=8'hd7;
        mem_19[14]=8'hab;
        mem_19[15]=8'h76;
        mem_19[16]=8'hca;
        mem_19[17]=8'h82;
        mem_19[18]=8'hc9;
        mem_19[19]=8'h7d;
        mem_19[20]=8'hfa;
        mem_19[21]=8'h59;
        mem_19[22]=8'h47;
        mem_19[23]=8'hf0;
        mem_19[24]=8'had;
        mem_19[25]=8'hd4;
        mem_19[26]=8'ha2;
        mem_19[27]=8'haf;
        mem_19[28]=8'h9c;
        mem_19[29]=8'ha4;
        mem_19[30]=8'h72;
        mem_19[31]=8'hc0;
        mem_19[32]=8'hb7;
        mem_19[33]=8'hfd;
        mem_19[34]=8'h93;
        mem_19[35]=8'h26;
        mem_19[36]=8'h36;
        mem_19[37]=8'h3f;
        mem_19[38]=8'hf7;
        mem_19[39]=8'hcc;
        mem_19[40]=8'h34;
        mem_19[41]=8'ha5;
        mem_19[42]=8'he5;
        mem_19[43]=8'hf1;
        mem_19[44]=8'h71;
        mem_19[45]=8'hd8;
        mem_19[46]=8'h31;
        mem_19[47]=8'h15;
        mem_19[48]=8'h4;
        mem_19[49]=8'hc7;
        mem_19[50]=8'h23;
        mem_19[51]=8'hc3;
        mem_19[52]=8'h18;
        mem_19[53]=8'h96;
        mem_19[54]=8'h5;
        mem_19[55]=8'h9a;
        mem_19[56]=8'h7;
        mem_19[57]=8'h12;
        mem_19[58]=8'h80;
        mem_19[59]=8'he2;
        mem_19[60]=8'heb;
        mem_19[61]=8'h27;
        mem_19[62]=8'hb2;
        mem_19[63]=8'h75;
        mem_19[64]=8'h9;
        mem_19[65]=8'h83;
        mem_19[66]=8'h2c;
        mem_19[67]=8'h1a;
        mem_19[68]=8'h1b;
        mem_19[69]=8'h6e;
        mem_19[70]=8'h5a;
        mem_19[71]=8'ha0;
        mem_19[72]=8'h52;
        mem_19[73]=8'h3b;
        mem_19[74]=8'hd6;
        mem_19[75]=8'hb3;
        mem_19[76]=8'h29;
        mem_19[77]=8'he3;
        mem_19[78]=8'h2f;
        mem_19[79]=8'h84;
        mem_19[80]=8'h53;
        mem_19[81]=8'hd1;
        mem_19[82]=8'h0;
        mem_19[83]=8'hed;
        mem_19[84]=8'h20;
        mem_19[85]=8'hfc;
        mem_19[86]=8'hb1;
        mem_19[87]=8'h5b;
        mem_19[88]=8'h6a;
        mem_19[89]=8'hcb;
        mem_19[90]=8'hbe;
        mem_19[91]=8'h39;
        mem_19[92]=8'h4a;
        mem_19[93]=8'h4c;
        mem_19[94]=8'h58;
        mem_19[95]=8'hcf;
        mem_19[96]=8'hd0;
        mem_19[97]=8'hef;
        mem_19[98]=8'haa;
        mem_19[99]=8'hfb;
        mem_19[100]=8'h43;
        mem_19[101]=8'h4d;
        mem_19[102]=8'h33;
        mem_19[103]=8'h85;
        mem_19[104]=8'h45;
        mem_19[105]=8'hf9;
        mem_19[106]=8'h2;
        mem_19[107]=8'h7f;
        mem_19[108]=8'h50;
        mem_19[109]=8'h3c;
        mem_19[110]=8'h9f;
        mem_19[111]=8'ha8;
        mem_19[112]=8'h51;
        mem_19[113]=8'ha3;
        mem_19[114]=8'h40;
        mem_19[115]=8'h8f;
        mem_19[116]=8'h92;
        mem_19[117]=8'h9d;
        mem_19[118]=8'h38;
        mem_19[119]=8'hf5;
        mem_19[120]=8'hbc;
        mem_19[121]=8'hb6;
        mem_19[122]=8'hda;
        mem_19[123]=8'h21;
        mem_19[124]=8'h10;
        mem_19[125]=8'hff;
        mem_19[126]=8'hf3;
        mem_19[127]=8'hd2;
        mem_19[128]=8'hcd;
        mem_19[129]=8'hc;
        mem_19[130]=8'h13;
        mem_19[131]=8'hec;
        mem_19[132]=8'h5f;
        mem_19[133]=8'h97;
        mem_19[134]=8'h44;
        mem_19[135]=8'h17;
        mem_19[136]=8'hc4;
        mem_19[137]=8'ha7;
        mem_19[138]=8'h7e;
        mem_19[139]=8'h3d;
        mem_19[140]=8'h64;
        mem_19[141]=8'h5d;
        mem_19[142]=8'h19;
        mem_19[143]=8'h73;
        mem_19[144]=8'h60;
        mem_19[145]=8'h81;
        mem_19[146]=8'h4f;
        mem_19[147]=8'hdc;
        mem_19[148]=8'h22;
        mem_19[149]=8'h2a;
        mem_19[150]=8'h90;
        mem_19[151]=8'h88;
        mem_19[152]=8'h46;
        mem_19[153]=8'hee;
        mem_19[154]=8'hb8;
        mem_19[155]=8'h14;
        mem_19[156]=8'hde;
        mem_19[157]=8'h5e;
        mem_19[158]=8'hb;
        mem_19[159]=8'hdb;
        mem_19[160]=8'he0;
        mem_19[161]=8'h32;
        mem_19[162]=8'h3a;
        mem_19[163]=8'ha;
        mem_19[164]=8'h49;
        mem_19[165]=8'h6;
        mem_19[166]=8'h24;
        mem_19[167]=8'h5c;
        mem_19[168]=8'hc2;
        mem_19[169]=8'hd3;
        mem_19[170]=8'hac;
        mem_19[171]=8'h62;
        mem_19[172]=8'h91;
        mem_19[173]=8'h95;
        mem_19[174]=8'he4;
        mem_19[175]=8'h79;
        mem_19[176]=8'he7;
        mem_19[177]=8'hc8;
        mem_19[178]=8'h37;
        mem_19[179]=8'h6d;
        mem_19[180]=8'h8d;
        mem_19[181]=8'hd5;
        mem_19[182]=8'h4e;
        mem_19[183]=8'ha9;
        mem_19[184]=8'h6c;
        mem_19[185]=8'h56;
        mem_19[186]=8'hf4;
        mem_19[187]=8'hea;
        mem_19[188]=8'h65;
        mem_19[189]=8'h7a;
        mem_19[190]=8'hae;
        mem_19[191]=8'h8;
        mem_19[192]=8'hba;
        mem_19[193]=8'h78;
        mem_19[194]=8'h25;
        mem_19[195]=8'h2e;
        mem_19[196]=8'h1c;
        mem_19[197]=8'ha6;
        mem_19[198]=8'hb4;
        mem_19[199]=8'hc6;
        mem_19[200]=8'he8;
        mem_19[201]=8'hdd;
        mem_19[202]=8'h74;
        mem_19[203]=8'h1f;
        mem_19[204]=8'h4b;
        mem_19[205]=8'hbd;
        mem_19[206]=8'h8b;
        mem_19[207]=8'h8a;
        mem_19[208]=8'h70;
        mem_19[209]=8'h3e;
        mem_19[210]=8'hb5;
        mem_19[211]=8'h66;
        mem_19[212]=8'h48;
        mem_19[213]=8'h3;
        mem_19[214]=8'hf6;
        mem_19[215]=8'he;
        mem_19[216]=8'h61;
        mem_19[217]=8'h35;
        mem_19[218]=8'h57;
        mem_19[219]=8'hb9;
        mem_19[220]=8'h86;
        mem_19[221]=8'hc1;
        mem_19[222]=8'h1d;
        mem_19[223]=8'h9e;
        mem_19[224]=8'he1;
        mem_19[225]=8'hf8;
        mem_19[226]=8'h98;
        mem_19[227]=8'h11;
        mem_19[228]=8'h69;
        mem_19[229]=8'hd9;
        mem_19[230]=8'h8e;
        mem_19[231]=8'h94;
        mem_19[232]=8'h9b;
        mem_19[233]=8'h1e;
        mem_19[234]=8'h87;
        mem_19[235]=8'he9;
        mem_19[236]=8'hce;
        mem_19[237]=8'h55;
        mem_19[238]=8'h28;
        mem_19[239]=8'hdf;
        mem_19[240]=8'h8c;
        mem_19[241]=8'ha1;
        mem_19[242]=8'h89;
        mem_19[243]=8'hd;
        mem_19[244]=8'hbf;
        mem_19[245]=8'he6;
        mem_19[246]=8'h42;
        mem_19[247]=8'h68;
        mem_19[248]=8'h41;
        mem_19[249]=8'h99;
        mem_19[250]=8'h2d;
        mem_19[251]=8'hf;
        mem_19[252]=8'hb0;
        mem_19[253]=8'h54;
        mem_19[254]=8'hbb;
        mem_19[255]=8'h16;
    end

    initial begin
        mem_20[0]=8'h63;
        mem_20[1]=8'h7c;
        mem_20[2]=8'h77;
        mem_20[3]=8'h7b;
        mem_20[4]=8'hf2;
        mem_20[5]=8'h6b;
        mem_20[6]=8'h6f;
        mem_20[7]=8'hc5;
        mem_20[8]=8'h30;
        mem_20[9]=8'h1;
        mem_20[10]=8'h67;
        mem_20[11]=8'h2b;
        mem_20[12]=8'hfe;
        mem_20[13]=8'hd7;
        mem_20[14]=8'hab;
        mem_20[15]=8'h76;
        mem_20[16]=8'hca;
        mem_20[17]=8'h82;
        mem_20[18]=8'hc9;
        mem_20[19]=8'h7d;
        mem_20[20]=8'hfa;
        mem_20[21]=8'h59;
        mem_20[22]=8'h47;
        mem_20[23]=8'hf0;
        mem_20[24]=8'had;
        mem_20[25]=8'hd4;
        mem_20[26]=8'ha2;
        mem_20[27]=8'haf;
        mem_20[28]=8'h9c;
        mem_20[29]=8'ha4;
        mem_20[30]=8'h72;
        mem_20[31]=8'hc0;
        mem_20[32]=8'hb7;
        mem_20[33]=8'hfd;
        mem_20[34]=8'h93;
        mem_20[35]=8'h26;
        mem_20[36]=8'h36;
        mem_20[37]=8'h3f;
        mem_20[38]=8'hf7;
        mem_20[39]=8'hcc;
        mem_20[40]=8'h34;
        mem_20[41]=8'ha5;
        mem_20[42]=8'he5;
        mem_20[43]=8'hf1;
        mem_20[44]=8'h71;
        mem_20[45]=8'hd8;
        mem_20[46]=8'h31;
        mem_20[47]=8'h15;
        mem_20[48]=8'h4;
        mem_20[49]=8'hc7;
        mem_20[50]=8'h23;
        mem_20[51]=8'hc3;
        mem_20[52]=8'h18;
        mem_20[53]=8'h96;
        mem_20[54]=8'h5;
        mem_20[55]=8'h9a;
        mem_20[56]=8'h7;
        mem_20[57]=8'h12;
        mem_20[58]=8'h80;
        mem_20[59]=8'he2;
        mem_20[60]=8'heb;
        mem_20[61]=8'h27;
        mem_20[62]=8'hb2;
        mem_20[63]=8'h75;
        mem_20[64]=8'h9;
        mem_20[65]=8'h83;
        mem_20[66]=8'h2c;
        mem_20[67]=8'h1a;
        mem_20[68]=8'h1b;
        mem_20[69]=8'h6e;
        mem_20[70]=8'h5a;
        mem_20[71]=8'ha0;
        mem_20[72]=8'h52;
        mem_20[73]=8'h3b;
        mem_20[74]=8'hd6;
        mem_20[75]=8'hb3;
        mem_20[76]=8'h29;
        mem_20[77]=8'he3;
        mem_20[78]=8'h2f;
        mem_20[79]=8'h84;
        mem_20[80]=8'h53;
        mem_20[81]=8'hd1;
        mem_20[82]=8'h0;
        mem_20[83]=8'hed;
        mem_20[84]=8'h20;
        mem_20[85]=8'hfc;
        mem_20[86]=8'hb1;
        mem_20[87]=8'h5b;
        mem_20[88]=8'h6a;
        mem_20[89]=8'hcb;
        mem_20[90]=8'hbe;
        mem_20[91]=8'h39;
        mem_20[92]=8'h4a;
        mem_20[93]=8'h4c;
        mem_20[94]=8'h58;
        mem_20[95]=8'hcf;
        mem_20[96]=8'hd0;
        mem_20[97]=8'hef;
        mem_20[98]=8'haa;
        mem_20[99]=8'hfb;
        mem_20[100]=8'h43;
        mem_20[101]=8'h4d;
        mem_20[102]=8'h33;
        mem_20[103]=8'h85;
        mem_20[104]=8'h45;
        mem_20[105]=8'hf9;
        mem_20[106]=8'h2;
        mem_20[107]=8'h7f;
        mem_20[108]=8'h50;
        mem_20[109]=8'h3c;
        mem_20[110]=8'h9f;
        mem_20[111]=8'ha8;
        mem_20[112]=8'h51;
        mem_20[113]=8'ha3;
        mem_20[114]=8'h40;
        mem_20[115]=8'h8f;
        mem_20[116]=8'h92;
        mem_20[117]=8'h9d;
        mem_20[118]=8'h38;
        mem_20[119]=8'hf5;
        mem_20[120]=8'hbc;
        mem_20[121]=8'hb6;
        mem_20[122]=8'hda;
        mem_20[123]=8'h21;
        mem_20[124]=8'h10;
        mem_20[125]=8'hff;
        mem_20[126]=8'hf3;
        mem_20[127]=8'hd2;
        mem_20[128]=8'hcd;
        mem_20[129]=8'hc;
        mem_20[130]=8'h13;
        mem_20[131]=8'hec;
        mem_20[132]=8'h5f;
        mem_20[133]=8'h97;
        mem_20[134]=8'h44;
        mem_20[135]=8'h17;
        mem_20[136]=8'hc4;
        mem_20[137]=8'ha7;
        mem_20[138]=8'h7e;
        mem_20[139]=8'h3d;
        mem_20[140]=8'h64;
        mem_20[141]=8'h5d;
        mem_20[142]=8'h19;
        mem_20[143]=8'h73;
        mem_20[144]=8'h60;
        mem_20[145]=8'h81;
        mem_20[146]=8'h4f;
        mem_20[147]=8'hdc;
        mem_20[148]=8'h22;
        mem_20[149]=8'h2a;
        mem_20[150]=8'h90;
        mem_20[151]=8'h88;
        mem_20[152]=8'h46;
        mem_20[153]=8'hee;
        mem_20[154]=8'hb8;
        mem_20[155]=8'h14;
        mem_20[156]=8'hde;
        mem_20[157]=8'h5e;
        mem_20[158]=8'hb;
        mem_20[159]=8'hdb;
        mem_20[160]=8'he0;
        mem_20[161]=8'h32;
        mem_20[162]=8'h3a;
        mem_20[163]=8'ha;
        mem_20[164]=8'h49;
        mem_20[165]=8'h6;
        mem_20[166]=8'h24;
        mem_20[167]=8'h5c;
        mem_20[168]=8'hc2;
        mem_20[169]=8'hd3;
        mem_20[170]=8'hac;
        mem_20[171]=8'h62;
        mem_20[172]=8'h91;
        mem_20[173]=8'h95;
        mem_20[174]=8'he4;
        mem_20[175]=8'h79;
        mem_20[176]=8'he7;
        mem_20[177]=8'hc8;
        mem_20[178]=8'h37;
        mem_20[179]=8'h6d;
        mem_20[180]=8'h8d;
        mem_20[181]=8'hd5;
        mem_20[182]=8'h4e;
        mem_20[183]=8'ha9;
        mem_20[184]=8'h6c;
        mem_20[185]=8'h56;
        mem_20[186]=8'hf4;
        mem_20[187]=8'hea;
        mem_20[188]=8'h65;
        mem_20[189]=8'h7a;
        mem_20[190]=8'hae;
        mem_20[191]=8'h8;
        mem_20[192]=8'hba;
        mem_20[193]=8'h78;
        mem_20[194]=8'h25;
        mem_20[195]=8'h2e;
        mem_20[196]=8'h1c;
        mem_20[197]=8'ha6;
        mem_20[198]=8'hb4;
        mem_20[199]=8'hc6;
        mem_20[200]=8'he8;
        mem_20[201]=8'hdd;
        mem_20[202]=8'h74;
        mem_20[203]=8'h1f;
        mem_20[204]=8'h4b;
        mem_20[205]=8'hbd;
        mem_20[206]=8'h8b;
        mem_20[207]=8'h8a;
        mem_20[208]=8'h70;
        mem_20[209]=8'h3e;
        mem_20[210]=8'hb5;
        mem_20[211]=8'h66;
        mem_20[212]=8'h48;
        mem_20[213]=8'h3;
        mem_20[214]=8'hf6;
        mem_20[215]=8'he;
        mem_20[216]=8'h61;
        mem_20[217]=8'h35;
        mem_20[218]=8'h57;
        mem_20[219]=8'hb9;
        mem_20[220]=8'h86;
        mem_20[221]=8'hc1;
        mem_20[222]=8'h1d;
        mem_20[223]=8'h9e;
        mem_20[224]=8'he1;
        mem_20[225]=8'hf8;
        mem_20[226]=8'h98;
        mem_20[227]=8'h11;
        mem_20[228]=8'h69;
        mem_20[229]=8'hd9;
        mem_20[230]=8'h8e;
        mem_20[231]=8'h94;
        mem_20[232]=8'h9b;
        mem_20[233]=8'h1e;
        mem_20[234]=8'h87;
        mem_20[235]=8'he9;
        mem_20[236]=8'hce;
        mem_20[237]=8'h55;
        mem_20[238]=8'h28;
        mem_20[239]=8'hdf;
        mem_20[240]=8'h8c;
        mem_20[241]=8'ha1;
        mem_20[242]=8'h89;
        mem_20[243]=8'hd;
        mem_20[244]=8'hbf;
        mem_20[245]=8'he6;
        mem_20[246]=8'h42;
        mem_20[247]=8'h68;
        mem_20[248]=8'h41;
        mem_20[249]=8'h99;
        mem_20[250]=8'h2d;
        mem_20[251]=8'hf;
        mem_20[252]=8'hb0;
        mem_20[253]=8'h54;
        mem_20[254]=8'hbb;
        mem_20[255]=8'h16;
    end

    initial begin
        mem_21[0]=8'h63;
        mem_21[1]=8'h7c;
        mem_21[2]=8'h77;
        mem_21[3]=8'h7b;
        mem_21[4]=8'hf2;
        mem_21[5]=8'h6b;
        mem_21[6]=8'h6f;
        mem_21[7]=8'hc5;
        mem_21[8]=8'h30;
        mem_21[9]=8'h1;
        mem_21[10]=8'h67;
        mem_21[11]=8'h2b;
        mem_21[12]=8'hfe;
        mem_21[13]=8'hd7;
        mem_21[14]=8'hab;
        mem_21[15]=8'h76;
        mem_21[16]=8'hca;
        mem_21[17]=8'h82;
        mem_21[18]=8'hc9;
        mem_21[19]=8'h7d;
        mem_21[20]=8'hfa;
        mem_21[21]=8'h59;
        mem_21[22]=8'h47;
        mem_21[23]=8'hf0;
        mem_21[24]=8'had;
        mem_21[25]=8'hd4;
        mem_21[26]=8'ha2;
        mem_21[27]=8'haf;
        mem_21[28]=8'h9c;
        mem_21[29]=8'ha4;
        mem_21[30]=8'h72;
        mem_21[31]=8'hc0;
        mem_21[32]=8'hb7;
        mem_21[33]=8'hfd;
        mem_21[34]=8'h93;
        mem_21[35]=8'h26;
        mem_21[36]=8'h36;
        mem_21[37]=8'h3f;
        mem_21[38]=8'hf7;
        mem_21[39]=8'hcc;
        mem_21[40]=8'h34;
        mem_21[41]=8'ha5;
        mem_21[42]=8'he5;
        mem_21[43]=8'hf1;
        mem_21[44]=8'h71;
        mem_21[45]=8'hd8;
        mem_21[46]=8'h31;
        mem_21[47]=8'h15;
        mem_21[48]=8'h4;
        mem_21[49]=8'hc7;
        mem_21[50]=8'h23;
        mem_21[51]=8'hc3;
        mem_21[52]=8'h18;
        mem_21[53]=8'h96;
        mem_21[54]=8'h5;
        mem_21[55]=8'h9a;
        mem_21[56]=8'h7;
        mem_21[57]=8'h12;
        mem_21[58]=8'h80;
        mem_21[59]=8'he2;
        mem_21[60]=8'heb;
        mem_21[61]=8'h27;
        mem_21[62]=8'hb2;
        mem_21[63]=8'h75;
        mem_21[64]=8'h9;
        mem_21[65]=8'h83;
        mem_21[66]=8'h2c;
        mem_21[67]=8'h1a;
        mem_21[68]=8'h1b;
        mem_21[69]=8'h6e;
        mem_21[70]=8'h5a;
        mem_21[71]=8'ha0;
        mem_21[72]=8'h52;
        mem_21[73]=8'h3b;
        mem_21[74]=8'hd6;
        mem_21[75]=8'hb3;
        mem_21[76]=8'h29;
        mem_21[77]=8'he3;
        mem_21[78]=8'h2f;
        mem_21[79]=8'h84;
        mem_21[80]=8'h53;
        mem_21[81]=8'hd1;
        mem_21[82]=8'h0;
        mem_21[83]=8'hed;
        mem_21[84]=8'h20;
        mem_21[85]=8'hfc;
        mem_21[86]=8'hb1;
        mem_21[87]=8'h5b;
        mem_21[88]=8'h6a;
        mem_21[89]=8'hcb;
        mem_21[90]=8'hbe;
        mem_21[91]=8'h39;
        mem_21[92]=8'h4a;
        mem_21[93]=8'h4c;
        mem_21[94]=8'h58;
        mem_21[95]=8'hcf;
        mem_21[96]=8'hd0;
        mem_21[97]=8'hef;
        mem_21[98]=8'haa;
        mem_21[99]=8'hfb;
        mem_21[100]=8'h43;
        mem_21[101]=8'h4d;
        mem_21[102]=8'h33;
        mem_21[103]=8'h85;
        mem_21[104]=8'h45;
        mem_21[105]=8'hf9;
        mem_21[106]=8'h2;
        mem_21[107]=8'h7f;
        mem_21[108]=8'h50;
        mem_21[109]=8'h3c;
        mem_21[110]=8'h9f;
        mem_21[111]=8'ha8;
        mem_21[112]=8'h51;
        mem_21[113]=8'ha3;
        mem_21[114]=8'h40;
        mem_21[115]=8'h8f;
        mem_21[116]=8'h92;
        mem_21[117]=8'h9d;
        mem_21[118]=8'h38;
        mem_21[119]=8'hf5;
        mem_21[120]=8'hbc;
        mem_21[121]=8'hb6;
        mem_21[122]=8'hda;
        mem_21[123]=8'h21;
        mem_21[124]=8'h10;
        mem_21[125]=8'hff;
        mem_21[126]=8'hf3;
        mem_21[127]=8'hd2;
        mem_21[128]=8'hcd;
        mem_21[129]=8'hc;
        mem_21[130]=8'h13;
        mem_21[131]=8'hec;
        mem_21[132]=8'h5f;
        mem_21[133]=8'h97;
        mem_21[134]=8'h44;
        mem_21[135]=8'h17;
        mem_21[136]=8'hc4;
        mem_21[137]=8'ha7;
        mem_21[138]=8'h7e;
        mem_21[139]=8'h3d;
        mem_21[140]=8'h64;
        mem_21[141]=8'h5d;
        mem_21[142]=8'h19;
        mem_21[143]=8'h73;
        mem_21[144]=8'h60;
        mem_21[145]=8'h81;
        mem_21[146]=8'h4f;
        mem_21[147]=8'hdc;
        mem_21[148]=8'h22;
        mem_21[149]=8'h2a;
        mem_21[150]=8'h90;
        mem_21[151]=8'h88;
        mem_21[152]=8'h46;
        mem_21[153]=8'hee;
        mem_21[154]=8'hb8;
        mem_21[155]=8'h14;
        mem_21[156]=8'hde;
        mem_21[157]=8'h5e;
        mem_21[158]=8'hb;
        mem_21[159]=8'hdb;
        mem_21[160]=8'he0;
        mem_21[161]=8'h32;
        mem_21[162]=8'h3a;
        mem_21[163]=8'ha;
        mem_21[164]=8'h49;
        mem_21[165]=8'h6;
        mem_21[166]=8'h24;
        mem_21[167]=8'h5c;
        mem_21[168]=8'hc2;
        mem_21[169]=8'hd3;
        mem_21[170]=8'hac;
        mem_21[171]=8'h62;
        mem_21[172]=8'h91;
        mem_21[173]=8'h95;
        mem_21[174]=8'he4;
        mem_21[175]=8'h79;
        mem_21[176]=8'he7;
        mem_21[177]=8'hc8;
        mem_21[178]=8'h37;
        mem_21[179]=8'h6d;
        mem_21[180]=8'h8d;
        mem_21[181]=8'hd5;
        mem_21[182]=8'h4e;
        mem_21[183]=8'ha9;
        mem_21[184]=8'h6c;
        mem_21[185]=8'h56;
        mem_21[186]=8'hf4;
        mem_21[187]=8'hea;
        mem_21[188]=8'h65;
        mem_21[189]=8'h7a;
        mem_21[190]=8'hae;
        mem_21[191]=8'h8;
        mem_21[192]=8'hba;
        mem_21[193]=8'h78;
        mem_21[194]=8'h25;
        mem_21[195]=8'h2e;
        mem_21[196]=8'h1c;
        mem_21[197]=8'ha6;
        mem_21[198]=8'hb4;
        mem_21[199]=8'hc6;
        mem_21[200]=8'he8;
        mem_21[201]=8'hdd;
        mem_21[202]=8'h74;
        mem_21[203]=8'h1f;
        mem_21[204]=8'h4b;
        mem_21[205]=8'hbd;
        mem_21[206]=8'h8b;
        mem_21[207]=8'h8a;
        mem_21[208]=8'h70;
        mem_21[209]=8'h3e;
        mem_21[210]=8'hb5;
        mem_21[211]=8'h66;
        mem_21[212]=8'h48;
        mem_21[213]=8'h3;
        mem_21[214]=8'hf6;
        mem_21[215]=8'he;
        mem_21[216]=8'h61;
        mem_21[217]=8'h35;
        mem_21[218]=8'h57;
        mem_21[219]=8'hb9;
        mem_21[220]=8'h86;
        mem_21[221]=8'hc1;
        mem_21[222]=8'h1d;
        mem_21[223]=8'h9e;
        mem_21[224]=8'he1;
        mem_21[225]=8'hf8;
        mem_21[226]=8'h98;
        mem_21[227]=8'h11;
        mem_21[228]=8'h69;
        mem_21[229]=8'hd9;
        mem_21[230]=8'h8e;
        mem_21[231]=8'h94;
        mem_21[232]=8'h9b;
        mem_21[233]=8'h1e;
        mem_21[234]=8'h87;
        mem_21[235]=8'he9;
        mem_21[236]=8'hce;
        mem_21[237]=8'h55;
        mem_21[238]=8'h28;
        mem_21[239]=8'hdf;
        mem_21[240]=8'h8c;
        mem_21[241]=8'ha1;
        mem_21[242]=8'h89;
        mem_21[243]=8'hd;
        mem_21[244]=8'hbf;
        mem_21[245]=8'he6;
        mem_21[246]=8'h42;
        mem_21[247]=8'h68;
        mem_21[248]=8'h41;
        mem_21[249]=8'h99;
        mem_21[250]=8'h2d;
        mem_21[251]=8'hf;
        mem_21[252]=8'hb0;
        mem_21[253]=8'h54;
        mem_21[254]=8'hbb;
        mem_21[255]=8'h16;
    end

    initial begin
        mem_22[0]=8'h63;
        mem_22[1]=8'h7c;
        mem_22[2]=8'h77;
        mem_22[3]=8'h7b;
        mem_22[4]=8'hf2;
        mem_22[5]=8'h6b;
        mem_22[6]=8'h6f;
        mem_22[7]=8'hc5;
        mem_22[8]=8'h30;
        mem_22[9]=8'h1;
        mem_22[10]=8'h67;
        mem_22[11]=8'h2b;
        mem_22[12]=8'hfe;
        mem_22[13]=8'hd7;
        mem_22[14]=8'hab;
        mem_22[15]=8'h76;
        mem_22[16]=8'hca;
        mem_22[17]=8'h82;
        mem_22[18]=8'hc9;
        mem_22[19]=8'h7d;
        mem_22[20]=8'hfa;
        mem_22[21]=8'h59;
        mem_22[22]=8'h47;
        mem_22[23]=8'hf0;
        mem_22[24]=8'had;
        mem_22[25]=8'hd4;
        mem_22[26]=8'ha2;
        mem_22[27]=8'haf;
        mem_22[28]=8'h9c;
        mem_22[29]=8'ha4;
        mem_22[30]=8'h72;
        mem_22[31]=8'hc0;
        mem_22[32]=8'hb7;
        mem_22[33]=8'hfd;
        mem_22[34]=8'h93;
        mem_22[35]=8'h26;
        mem_22[36]=8'h36;
        mem_22[37]=8'h3f;
        mem_22[38]=8'hf7;
        mem_22[39]=8'hcc;
        mem_22[40]=8'h34;
        mem_22[41]=8'ha5;
        mem_22[42]=8'he5;
        mem_22[43]=8'hf1;
        mem_22[44]=8'h71;
        mem_22[45]=8'hd8;
        mem_22[46]=8'h31;
        mem_22[47]=8'h15;
        mem_22[48]=8'h4;
        mem_22[49]=8'hc7;
        mem_22[50]=8'h23;
        mem_22[51]=8'hc3;
        mem_22[52]=8'h18;
        mem_22[53]=8'h96;
        mem_22[54]=8'h5;
        mem_22[55]=8'h9a;
        mem_22[56]=8'h7;
        mem_22[57]=8'h12;
        mem_22[58]=8'h80;
        mem_22[59]=8'he2;
        mem_22[60]=8'heb;
        mem_22[61]=8'h27;
        mem_22[62]=8'hb2;
        mem_22[63]=8'h75;
        mem_22[64]=8'h9;
        mem_22[65]=8'h83;
        mem_22[66]=8'h2c;
        mem_22[67]=8'h1a;
        mem_22[68]=8'h1b;
        mem_22[69]=8'h6e;
        mem_22[70]=8'h5a;
        mem_22[71]=8'ha0;
        mem_22[72]=8'h52;
        mem_22[73]=8'h3b;
        mem_22[74]=8'hd6;
        mem_22[75]=8'hb3;
        mem_22[76]=8'h29;
        mem_22[77]=8'he3;
        mem_22[78]=8'h2f;
        mem_22[79]=8'h84;
        mem_22[80]=8'h53;
        mem_22[81]=8'hd1;
        mem_22[82]=8'h0;
        mem_22[83]=8'hed;
        mem_22[84]=8'h20;
        mem_22[85]=8'hfc;
        mem_22[86]=8'hb1;
        mem_22[87]=8'h5b;
        mem_22[88]=8'h6a;
        mem_22[89]=8'hcb;
        mem_22[90]=8'hbe;
        mem_22[91]=8'h39;
        mem_22[92]=8'h4a;
        mem_22[93]=8'h4c;
        mem_22[94]=8'h58;
        mem_22[95]=8'hcf;
        mem_22[96]=8'hd0;
        mem_22[97]=8'hef;
        mem_22[98]=8'haa;
        mem_22[99]=8'hfb;
        mem_22[100]=8'h43;
        mem_22[101]=8'h4d;
        mem_22[102]=8'h33;
        mem_22[103]=8'h85;
        mem_22[104]=8'h45;
        mem_22[105]=8'hf9;
        mem_22[106]=8'h2;
        mem_22[107]=8'h7f;
        mem_22[108]=8'h50;
        mem_22[109]=8'h3c;
        mem_22[110]=8'h9f;
        mem_22[111]=8'ha8;
        mem_22[112]=8'h51;
        mem_22[113]=8'ha3;
        mem_22[114]=8'h40;
        mem_22[115]=8'h8f;
        mem_22[116]=8'h92;
        mem_22[117]=8'h9d;
        mem_22[118]=8'h38;
        mem_22[119]=8'hf5;
        mem_22[120]=8'hbc;
        mem_22[121]=8'hb6;
        mem_22[122]=8'hda;
        mem_22[123]=8'h21;
        mem_22[124]=8'h10;
        mem_22[125]=8'hff;
        mem_22[126]=8'hf3;
        mem_22[127]=8'hd2;
        mem_22[128]=8'hcd;
        mem_22[129]=8'hc;
        mem_22[130]=8'h13;
        mem_22[131]=8'hec;
        mem_22[132]=8'h5f;
        mem_22[133]=8'h97;
        mem_22[134]=8'h44;
        mem_22[135]=8'h17;
        mem_22[136]=8'hc4;
        mem_22[137]=8'ha7;
        mem_22[138]=8'h7e;
        mem_22[139]=8'h3d;
        mem_22[140]=8'h64;
        mem_22[141]=8'h5d;
        mem_22[142]=8'h19;
        mem_22[143]=8'h73;
        mem_22[144]=8'h60;
        mem_22[145]=8'h81;
        mem_22[146]=8'h4f;
        mem_22[147]=8'hdc;
        mem_22[148]=8'h22;
        mem_22[149]=8'h2a;
        mem_22[150]=8'h90;
        mem_22[151]=8'h88;
        mem_22[152]=8'h46;
        mem_22[153]=8'hee;
        mem_22[154]=8'hb8;
        mem_22[155]=8'h14;
        mem_22[156]=8'hde;
        mem_22[157]=8'h5e;
        mem_22[158]=8'hb;
        mem_22[159]=8'hdb;
        mem_22[160]=8'he0;
        mem_22[161]=8'h32;
        mem_22[162]=8'h3a;
        mem_22[163]=8'ha;
        mem_22[164]=8'h49;
        mem_22[165]=8'h6;
        mem_22[166]=8'h24;
        mem_22[167]=8'h5c;
        mem_22[168]=8'hc2;
        mem_22[169]=8'hd3;
        mem_22[170]=8'hac;
        mem_22[171]=8'h62;
        mem_22[172]=8'h91;
        mem_22[173]=8'h95;
        mem_22[174]=8'he4;
        mem_22[175]=8'h79;
        mem_22[176]=8'he7;
        mem_22[177]=8'hc8;
        mem_22[178]=8'h37;
        mem_22[179]=8'h6d;
        mem_22[180]=8'h8d;
        mem_22[181]=8'hd5;
        mem_22[182]=8'h4e;
        mem_22[183]=8'ha9;
        mem_22[184]=8'h6c;
        mem_22[185]=8'h56;
        mem_22[186]=8'hf4;
        mem_22[187]=8'hea;
        mem_22[188]=8'h65;
        mem_22[189]=8'h7a;
        mem_22[190]=8'hae;
        mem_22[191]=8'h8;
        mem_22[192]=8'hba;
        mem_22[193]=8'h78;
        mem_22[194]=8'h25;
        mem_22[195]=8'h2e;
        mem_22[196]=8'h1c;
        mem_22[197]=8'ha6;
        mem_22[198]=8'hb4;
        mem_22[199]=8'hc6;
        mem_22[200]=8'he8;
        mem_22[201]=8'hdd;
        mem_22[202]=8'h74;
        mem_22[203]=8'h1f;
        mem_22[204]=8'h4b;
        mem_22[205]=8'hbd;
        mem_22[206]=8'h8b;
        mem_22[207]=8'h8a;
        mem_22[208]=8'h70;
        mem_22[209]=8'h3e;
        mem_22[210]=8'hb5;
        mem_22[211]=8'h66;
        mem_22[212]=8'h48;
        mem_22[213]=8'h3;
        mem_22[214]=8'hf6;
        mem_22[215]=8'he;
        mem_22[216]=8'h61;
        mem_22[217]=8'h35;
        mem_22[218]=8'h57;
        mem_22[219]=8'hb9;
        mem_22[220]=8'h86;
        mem_22[221]=8'hc1;
        mem_22[222]=8'h1d;
        mem_22[223]=8'h9e;
        mem_22[224]=8'he1;
        mem_22[225]=8'hf8;
        mem_22[226]=8'h98;
        mem_22[227]=8'h11;
        mem_22[228]=8'h69;
        mem_22[229]=8'hd9;
        mem_22[230]=8'h8e;
        mem_22[231]=8'h94;
        mem_22[232]=8'h9b;
        mem_22[233]=8'h1e;
        mem_22[234]=8'h87;
        mem_22[235]=8'he9;
        mem_22[236]=8'hce;
        mem_22[237]=8'h55;
        mem_22[238]=8'h28;
        mem_22[239]=8'hdf;
        mem_22[240]=8'h8c;
        mem_22[241]=8'ha1;
        mem_22[242]=8'h89;
        mem_22[243]=8'hd;
        mem_22[244]=8'hbf;
        mem_22[245]=8'he6;
        mem_22[246]=8'h42;
        mem_22[247]=8'h68;
        mem_22[248]=8'h41;
        mem_22[249]=8'h99;
        mem_22[250]=8'h2d;
        mem_22[251]=8'hf;
        mem_22[252]=8'hb0;
        mem_22[253]=8'h54;
        mem_22[254]=8'hbb;
        mem_22[255]=8'h16;
    end

    initial begin
        mem_23[0]=8'h63;
        mem_23[1]=8'h7c;
        mem_23[2]=8'h77;
        mem_23[3]=8'h7b;
        mem_23[4]=8'hf2;
        mem_23[5]=8'h6b;
        mem_23[6]=8'h6f;
        mem_23[7]=8'hc5;
        mem_23[8]=8'h30;
        mem_23[9]=8'h1;
        mem_23[10]=8'h67;
        mem_23[11]=8'h2b;
        mem_23[12]=8'hfe;
        mem_23[13]=8'hd7;
        mem_23[14]=8'hab;
        mem_23[15]=8'h76;
        mem_23[16]=8'hca;
        mem_23[17]=8'h82;
        mem_23[18]=8'hc9;
        mem_23[19]=8'h7d;
        mem_23[20]=8'hfa;
        mem_23[21]=8'h59;
        mem_23[22]=8'h47;
        mem_23[23]=8'hf0;
        mem_23[24]=8'had;
        mem_23[25]=8'hd4;
        mem_23[26]=8'ha2;
        mem_23[27]=8'haf;
        mem_23[28]=8'h9c;
        mem_23[29]=8'ha4;
        mem_23[30]=8'h72;
        mem_23[31]=8'hc0;
        mem_23[32]=8'hb7;
        mem_23[33]=8'hfd;
        mem_23[34]=8'h93;
        mem_23[35]=8'h26;
        mem_23[36]=8'h36;
        mem_23[37]=8'h3f;
        mem_23[38]=8'hf7;
        mem_23[39]=8'hcc;
        mem_23[40]=8'h34;
        mem_23[41]=8'ha5;
        mem_23[42]=8'he5;
        mem_23[43]=8'hf1;
        mem_23[44]=8'h71;
        mem_23[45]=8'hd8;
        mem_23[46]=8'h31;
        mem_23[47]=8'h15;
        mem_23[48]=8'h4;
        mem_23[49]=8'hc7;
        mem_23[50]=8'h23;
        mem_23[51]=8'hc3;
        mem_23[52]=8'h18;
        mem_23[53]=8'h96;
        mem_23[54]=8'h5;
        mem_23[55]=8'h9a;
        mem_23[56]=8'h7;
        mem_23[57]=8'h12;
        mem_23[58]=8'h80;
        mem_23[59]=8'he2;
        mem_23[60]=8'heb;
        mem_23[61]=8'h27;
        mem_23[62]=8'hb2;
        mem_23[63]=8'h75;
        mem_23[64]=8'h9;
        mem_23[65]=8'h83;
        mem_23[66]=8'h2c;
        mem_23[67]=8'h1a;
        mem_23[68]=8'h1b;
        mem_23[69]=8'h6e;
        mem_23[70]=8'h5a;
        mem_23[71]=8'ha0;
        mem_23[72]=8'h52;
        mem_23[73]=8'h3b;
        mem_23[74]=8'hd6;
        mem_23[75]=8'hb3;
        mem_23[76]=8'h29;
        mem_23[77]=8'he3;
        mem_23[78]=8'h2f;
        mem_23[79]=8'h84;
        mem_23[80]=8'h53;
        mem_23[81]=8'hd1;
        mem_23[82]=8'h0;
        mem_23[83]=8'hed;
        mem_23[84]=8'h20;
        mem_23[85]=8'hfc;
        mem_23[86]=8'hb1;
        mem_23[87]=8'h5b;
        mem_23[88]=8'h6a;
        mem_23[89]=8'hcb;
        mem_23[90]=8'hbe;
        mem_23[91]=8'h39;
        mem_23[92]=8'h4a;
        mem_23[93]=8'h4c;
        mem_23[94]=8'h58;
        mem_23[95]=8'hcf;
        mem_23[96]=8'hd0;
        mem_23[97]=8'hef;
        mem_23[98]=8'haa;
        mem_23[99]=8'hfb;
        mem_23[100]=8'h43;
        mem_23[101]=8'h4d;
        mem_23[102]=8'h33;
        mem_23[103]=8'h85;
        mem_23[104]=8'h45;
        mem_23[105]=8'hf9;
        mem_23[106]=8'h2;
        mem_23[107]=8'h7f;
        mem_23[108]=8'h50;
        mem_23[109]=8'h3c;
        mem_23[110]=8'h9f;
        mem_23[111]=8'ha8;
        mem_23[112]=8'h51;
        mem_23[113]=8'ha3;
        mem_23[114]=8'h40;
        mem_23[115]=8'h8f;
        mem_23[116]=8'h92;
        mem_23[117]=8'h9d;
        mem_23[118]=8'h38;
        mem_23[119]=8'hf5;
        mem_23[120]=8'hbc;
        mem_23[121]=8'hb6;
        mem_23[122]=8'hda;
        mem_23[123]=8'h21;
        mem_23[124]=8'h10;
        mem_23[125]=8'hff;
        mem_23[126]=8'hf3;
        mem_23[127]=8'hd2;
        mem_23[128]=8'hcd;
        mem_23[129]=8'hc;
        mem_23[130]=8'h13;
        mem_23[131]=8'hec;
        mem_23[132]=8'h5f;
        mem_23[133]=8'h97;
        mem_23[134]=8'h44;
        mem_23[135]=8'h17;
        mem_23[136]=8'hc4;
        mem_23[137]=8'ha7;
        mem_23[138]=8'h7e;
        mem_23[139]=8'h3d;
        mem_23[140]=8'h64;
        mem_23[141]=8'h5d;
        mem_23[142]=8'h19;
        mem_23[143]=8'h73;
        mem_23[144]=8'h60;
        mem_23[145]=8'h81;
        mem_23[146]=8'h4f;
        mem_23[147]=8'hdc;
        mem_23[148]=8'h22;
        mem_23[149]=8'h2a;
        mem_23[150]=8'h90;
        mem_23[151]=8'h88;
        mem_23[152]=8'h46;
        mem_23[153]=8'hee;
        mem_23[154]=8'hb8;
        mem_23[155]=8'h14;
        mem_23[156]=8'hde;
        mem_23[157]=8'h5e;
        mem_23[158]=8'hb;
        mem_23[159]=8'hdb;
        mem_23[160]=8'he0;
        mem_23[161]=8'h32;
        mem_23[162]=8'h3a;
        mem_23[163]=8'ha;
        mem_23[164]=8'h49;
        mem_23[165]=8'h6;
        mem_23[166]=8'h24;
        mem_23[167]=8'h5c;
        mem_23[168]=8'hc2;
        mem_23[169]=8'hd3;
        mem_23[170]=8'hac;
        mem_23[171]=8'h62;
        mem_23[172]=8'h91;
        mem_23[173]=8'h95;
        mem_23[174]=8'he4;
        mem_23[175]=8'h79;
        mem_23[176]=8'he7;
        mem_23[177]=8'hc8;
        mem_23[178]=8'h37;
        mem_23[179]=8'h6d;
        mem_23[180]=8'h8d;
        mem_23[181]=8'hd5;
        mem_23[182]=8'h4e;
        mem_23[183]=8'ha9;
        mem_23[184]=8'h6c;
        mem_23[185]=8'h56;
        mem_23[186]=8'hf4;
        mem_23[187]=8'hea;
        mem_23[188]=8'h65;
        mem_23[189]=8'h7a;
        mem_23[190]=8'hae;
        mem_23[191]=8'h8;
        mem_23[192]=8'hba;
        mem_23[193]=8'h78;
        mem_23[194]=8'h25;
        mem_23[195]=8'h2e;
        mem_23[196]=8'h1c;
        mem_23[197]=8'ha6;
        mem_23[198]=8'hb4;
        mem_23[199]=8'hc6;
        mem_23[200]=8'he8;
        mem_23[201]=8'hdd;
        mem_23[202]=8'h74;
        mem_23[203]=8'h1f;
        mem_23[204]=8'h4b;
        mem_23[205]=8'hbd;
        mem_23[206]=8'h8b;
        mem_23[207]=8'h8a;
        mem_23[208]=8'h70;
        mem_23[209]=8'h3e;
        mem_23[210]=8'hb5;
        mem_23[211]=8'h66;
        mem_23[212]=8'h48;
        mem_23[213]=8'h3;
        mem_23[214]=8'hf6;
        mem_23[215]=8'he;
        mem_23[216]=8'h61;
        mem_23[217]=8'h35;
        mem_23[218]=8'h57;
        mem_23[219]=8'hb9;
        mem_23[220]=8'h86;
        mem_23[221]=8'hc1;
        mem_23[222]=8'h1d;
        mem_23[223]=8'h9e;
        mem_23[224]=8'he1;
        mem_23[225]=8'hf8;
        mem_23[226]=8'h98;
        mem_23[227]=8'h11;
        mem_23[228]=8'h69;
        mem_23[229]=8'hd9;
        mem_23[230]=8'h8e;
        mem_23[231]=8'h94;
        mem_23[232]=8'h9b;
        mem_23[233]=8'h1e;
        mem_23[234]=8'h87;
        mem_23[235]=8'he9;
        mem_23[236]=8'hce;
        mem_23[237]=8'h55;
        mem_23[238]=8'h28;
        mem_23[239]=8'hdf;
        mem_23[240]=8'h8c;
        mem_23[241]=8'ha1;
        mem_23[242]=8'h89;
        mem_23[243]=8'hd;
        mem_23[244]=8'hbf;
        mem_23[245]=8'he6;
        mem_23[246]=8'h42;
        mem_23[247]=8'h68;
        mem_23[248]=8'h41;
        mem_23[249]=8'h99;
        mem_23[250]=8'h2d;
        mem_23[251]=8'hf;
        mem_23[252]=8'hb0;
        mem_23[253]=8'h54;
        mem_23[254]=8'hbb;
        mem_23[255]=8'h16;
    end

    initial begin
        mem_24[0]=8'h0;
        mem_24[1]=8'h2;
        mem_24[2]=8'h4;
        mem_24[3]=8'h6;
        mem_24[4]=8'h8;
        mem_24[5]=8'ha;
        mem_24[6]=8'hc;
        mem_24[7]=8'he;
        mem_24[8]=8'h10;
        mem_24[9]=8'h12;
        mem_24[10]=8'h14;
        mem_24[11]=8'h16;
        mem_24[12]=8'h18;
        mem_24[13]=8'h1a;
        mem_24[14]=8'h1c;
        mem_24[15]=8'h1e;
        mem_24[16]=8'h20;
        mem_24[17]=8'h22;
        mem_24[18]=8'h24;
        mem_24[19]=8'h26;
        mem_24[20]=8'h28;
        mem_24[21]=8'h2a;
        mem_24[22]=8'h2c;
        mem_24[23]=8'h2e;
        mem_24[24]=8'h30;
        mem_24[25]=8'h32;
        mem_24[26]=8'h34;
        mem_24[27]=8'h36;
        mem_24[28]=8'h38;
        mem_24[29]=8'h3a;
        mem_24[30]=8'h3c;
        mem_24[31]=8'h3e;
        mem_24[32]=8'h40;
        mem_24[33]=8'h42;
        mem_24[34]=8'h44;
        mem_24[35]=8'h46;
        mem_24[36]=8'h48;
        mem_24[37]=8'h4a;
        mem_24[38]=8'h4c;
        mem_24[39]=8'h4e;
        mem_24[40]=8'h50;
        mem_24[41]=8'h52;
        mem_24[42]=8'h54;
        mem_24[43]=8'h56;
        mem_24[44]=8'h58;
        mem_24[45]=8'h5a;
        mem_24[46]=8'h5c;
        mem_24[47]=8'h5e;
        mem_24[48]=8'h60;
        mem_24[49]=8'h62;
        mem_24[50]=8'h64;
        mem_24[51]=8'h66;
        mem_24[52]=8'h68;
        mem_24[53]=8'h6a;
        mem_24[54]=8'h6c;
        mem_24[55]=8'h6e;
        mem_24[56]=8'h70;
        mem_24[57]=8'h72;
        mem_24[58]=8'h74;
        mem_24[59]=8'h76;
        mem_24[60]=8'h78;
        mem_24[61]=8'h7a;
        mem_24[62]=8'h7c;
        mem_24[63]=8'h7e;
        mem_24[64]=8'h80;
        mem_24[65]=8'h82;
        mem_24[66]=8'h84;
        mem_24[67]=8'h86;
        mem_24[68]=8'h88;
        mem_24[69]=8'h8a;
        mem_24[70]=8'h8c;
        mem_24[71]=8'h8e;
        mem_24[72]=8'h90;
        mem_24[73]=8'h92;
        mem_24[74]=8'h94;
        mem_24[75]=8'h96;
        mem_24[76]=8'h98;
        mem_24[77]=8'h9a;
        mem_24[78]=8'h9c;
        mem_24[79]=8'h9e;
        mem_24[80]=8'ha0;
        mem_24[81]=8'ha2;
        mem_24[82]=8'ha4;
        mem_24[83]=8'ha6;
        mem_24[84]=8'ha8;
        mem_24[85]=8'haa;
        mem_24[86]=8'hac;
        mem_24[87]=8'hae;
        mem_24[88]=8'hb0;
        mem_24[89]=8'hb2;
        mem_24[90]=8'hb4;
        mem_24[91]=8'hb6;
        mem_24[92]=8'hb8;
        mem_24[93]=8'hba;
        mem_24[94]=8'hbc;
        mem_24[95]=8'hbe;
        mem_24[96]=8'hc0;
        mem_24[97]=8'hc2;
        mem_24[98]=8'hc4;
        mem_24[99]=8'hc6;
        mem_24[100]=8'hc8;
        mem_24[101]=8'hca;
        mem_24[102]=8'hcc;
        mem_24[103]=8'hce;
        mem_24[104]=8'hd0;
        mem_24[105]=8'hd2;
        mem_24[106]=8'hd4;
        mem_24[107]=8'hd6;
        mem_24[108]=8'hd8;
        mem_24[109]=8'hda;
        mem_24[110]=8'hdc;
        mem_24[111]=8'hde;
        mem_24[112]=8'he0;
        mem_24[113]=8'he2;
        mem_24[114]=8'he4;
        mem_24[115]=8'he6;
        mem_24[116]=8'he8;
        mem_24[117]=8'hea;
        mem_24[118]=8'hec;
        mem_24[119]=8'hee;
        mem_24[120]=8'hf0;
        mem_24[121]=8'hf2;
        mem_24[122]=8'hf4;
        mem_24[123]=8'hf6;
        mem_24[124]=8'hf8;
        mem_24[125]=8'hfa;
        mem_24[126]=8'hfc;
        mem_24[127]=8'hfe;
        mem_24[128]=8'h1b;
        mem_24[129]=8'h19;
        mem_24[130]=8'h1f;
        mem_24[131]=8'h1d;
        mem_24[132]=8'h13;
        mem_24[133]=8'h11;
        mem_24[134]=8'h17;
        mem_24[135]=8'h15;
        mem_24[136]=8'hb;
        mem_24[137]=8'h9;
        mem_24[138]=8'hf;
        mem_24[139]=8'hd;
        mem_24[140]=8'h3;
        mem_24[141]=8'h1;
        mem_24[142]=8'h7;
        mem_24[143]=8'h5;
        mem_24[144]=8'h3b;
        mem_24[145]=8'h39;
        mem_24[146]=8'h3f;
        mem_24[147]=8'h3d;
        mem_24[148]=8'h33;
        mem_24[149]=8'h31;
        mem_24[150]=8'h37;
        mem_24[151]=8'h35;
        mem_24[152]=8'h2b;
        mem_24[153]=8'h29;
        mem_24[154]=8'h2f;
        mem_24[155]=8'h2d;
        mem_24[156]=8'h23;
        mem_24[157]=8'h21;
        mem_24[158]=8'h27;
        mem_24[159]=8'h25;
        mem_24[160]=8'h5b;
        mem_24[161]=8'h59;
        mem_24[162]=8'h5f;
        mem_24[163]=8'h5d;
        mem_24[164]=8'h53;
        mem_24[165]=8'h51;
        mem_24[166]=8'h57;
        mem_24[167]=8'h55;
        mem_24[168]=8'h4b;
        mem_24[169]=8'h49;
        mem_24[170]=8'h4f;
        mem_24[171]=8'h4d;
        mem_24[172]=8'h43;
        mem_24[173]=8'h41;
        mem_24[174]=8'h47;
        mem_24[175]=8'h45;
        mem_24[176]=8'h7b;
        mem_24[177]=8'h79;
        mem_24[178]=8'h7f;
        mem_24[179]=8'h7d;
        mem_24[180]=8'h73;
        mem_24[181]=8'h71;
        mem_24[182]=8'h77;
        mem_24[183]=8'h75;
        mem_24[184]=8'h6b;
        mem_24[185]=8'h69;
        mem_24[186]=8'h6f;
        mem_24[187]=8'h6d;
        mem_24[188]=8'h63;
        mem_24[189]=8'h61;
        mem_24[190]=8'h67;
        mem_24[191]=8'h65;
        mem_24[192]=8'h9b;
        mem_24[193]=8'h99;
        mem_24[194]=8'h9f;
        mem_24[195]=8'h9d;
        mem_24[196]=8'h93;
        mem_24[197]=8'h91;
        mem_24[198]=8'h97;
        mem_24[199]=8'h95;
        mem_24[200]=8'h8b;
        mem_24[201]=8'h89;
        mem_24[202]=8'h8f;
        mem_24[203]=8'h8d;
        mem_24[204]=8'h83;
        mem_24[205]=8'h81;
        mem_24[206]=8'h87;
        mem_24[207]=8'h85;
        mem_24[208]=8'hbb;
        mem_24[209]=8'hb9;
        mem_24[210]=8'hbf;
        mem_24[211]=8'hbd;
        mem_24[212]=8'hb3;
        mem_24[213]=8'hb1;
        mem_24[214]=8'hb7;
        mem_24[215]=8'hb5;
        mem_24[216]=8'hab;
        mem_24[217]=8'ha9;
        mem_24[218]=8'haf;
        mem_24[219]=8'had;
        mem_24[220]=8'ha3;
        mem_24[221]=8'ha1;
        mem_24[222]=8'ha7;
        mem_24[223]=8'ha5;
        mem_24[224]=8'hdb;
        mem_24[225]=8'hd9;
        mem_24[226]=8'hdf;
        mem_24[227]=8'hdd;
        mem_24[228]=8'hd3;
        mem_24[229]=8'hd1;
        mem_24[230]=8'hd7;
        mem_24[231]=8'hd5;
        mem_24[232]=8'hcb;
        mem_24[233]=8'hc9;
        mem_24[234]=8'hcf;
        mem_24[235]=8'hcd;
        mem_24[236]=8'hc3;
        mem_24[237]=8'hc1;
        mem_24[238]=8'hc7;
        mem_24[239]=8'hc5;
        mem_24[240]=8'hfb;
        mem_24[241]=8'hf9;
        mem_24[242]=8'hff;
        mem_24[243]=8'hfd;
        mem_24[244]=8'hf3;
        mem_24[245]=8'hf1;
        mem_24[246]=8'hf7;
        mem_24[247]=8'hf5;
        mem_24[248]=8'heb;
        mem_24[249]=8'he9;
        mem_24[250]=8'hef;
        mem_24[251]=8'hed;
        mem_24[252]=8'he3;
        mem_24[253]=8'he1;
        mem_24[254]=8'he7;
        mem_24[255]=8'he5;
    end

    initial begin
        mem_25[0]=8'h0;
        mem_25[1]=8'h3;
        mem_25[2]=8'h6;
        mem_25[3]=8'h5;
        mem_25[4]=8'hc;
        mem_25[5]=8'hf;
        mem_25[6]=8'ha;
        mem_25[7]=8'h9;
        mem_25[8]=8'h18;
        mem_25[9]=8'h1b;
        mem_25[10]=8'h1e;
        mem_25[11]=8'h1d;
        mem_25[12]=8'h14;
        mem_25[13]=8'h17;
        mem_25[14]=8'h12;
        mem_25[15]=8'h11;
        mem_25[16]=8'h30;
        mem_25[17]=8'h33;
        mem_25[18]=8'h36;
        mem_25[19]=8'h35;
        mem_25[20]=8'h3c;
        mem_25[21]=8'h3f;
        mem_25[22]=8'h3a;
        mem_25[23]=8'h39;
        mem_25[24]=8'h28;
        mem_25[25]=8'h2b;
        mem_25[26]=8'h2e;
        mem_25[27]=8'h2d;
        mem_25[28]=8'h24;
        mem_25[29]=8'h27;
        mem_25[30]=8'h22;
        mem_25[31]=8'h21;
        mem_25[32]=8'h60;
        mem_25[33]=8'h63;
        mem_25[34]=8'h66;
        mem_25[35]=8'h65;
        mem_25[36]=8'h6c;
        mem_25[37]=8'h6f;
        mem_25[38]=8'h6a;
        mem_25[39]=8'h69;
        mem_25[40]=8'h78;
        mem_25[41]=8'h7b;
        mem_25[42]=8'h7e;
        mem_25[43]=8'h7d;
        mem_25[44]=8'h74;
        mem_25[45]=8'h77;
        mem_25[46]=8'h72;
        mem_25[47]=8'h71;
        mem_25[48]=8'h50;
        mem_25[49]=8'h53;
        mem_25[50]=8'h56;
        mem_25[51]=8'h55;
        mem_25[52]=8'h5c;
        mem_25[53]=8'h5f;
        mem_25[54]=8'h5a;
        mem_25[55]=8'h59;
        mem_25[56]=8'h48;
        mem_25[57]=8'h4b;
        mem_25[58]=8'h4e;
        mem_25[59]=8'h4d;
        mem_25[60]=8'h44;
        mem_25[61]=8'h47;
        mem_25[62]=8'h42;
        mem_25[63]=8'h41;
        mem_25[64]=8'hc0;
        mem_25[65]=8'hc3;
        mem_25[66]=8'hc6;
        mem_25[67]=8'hc5;
        mem_25[68]=8'hcc;
        mem_25[69]=8'hcf;
        mem_25[70]=8'hca;
        mem_25[71]=8'hc9;
        mem_25[72]=8'hd8;
        mem_25[73]=8'hdb;
        mem_25[74]=8'hde;
        mem_25[75]=8'hdd;
        mem_25[76]=8'hd4;
        mem_25[77]=8'hd7;
        mem_25[78]=8'hd2;
        mem_25[79]=8'hd1;
        mem_25[80]=8'hf0;
        mem_25[81]=8'hf3;
        mem_25[82]=8'hf6;
        mem_25[83]=8'hf5;
        mem_25[84]=8'hfc;
        mem_25[85]=8'hff;
        mem_25[86]=8'hfa;
        mem_25[87]=8'hf9;
        mem_25[88]=8'he8;
        mem_25[89]=8'heb;
        mem_25[90]=8'hee;
        mem_25[91]=8'hed;
        mem_25[92]=8'he4;
        mem_25[93]=8'he7;
        mem_25[94]=8'he2;
        mem_25[95]=8'he1;
        mem_25[96]=8'ha0;
        mem_25[97]=8'ha3;
        mem_25[98]=8'ha6;
        mem_25[99]=8'ha5;
        mem_25[100]=8'hac;
        mem_25[101]=8'haf;
        mem_25[102]=8'haa;
        mem_25[103]=8'ha9;
        mem_25[104]=8'hb8;
        mem_25[105]=8'hbb;
        mem_25[106]=8'hbe;
        mem_25[107]=8'hbd;
        mem_25[108]=8'hb4;
        mem_25[109]=8'hb7;
        mem_25[110]=8'hb2;
        mem_25[111]=8'hb1;
        mem_25[112]=8'h90;
        mem_25[113]=8'h93;
        mem_25[114]=8'h96;
        mem_25[115]=8'h95;
        mem_25[116]=8'h9c;
        mem_25[117]=8'h9f;
        mem_25[118]=8'h9a;
        mem_25[119]=8'h99;
        mem_25[120]=8'h88;
        mem_25[121]=8'h8b;
        mem_25[122]=8'h8e;
        mem_25[123]=8'h8d;
        mem_25[124]=8'h84;
        mem_25[125]=8'h87;
        mem_25[126]=8'h82;
        mem_25[127]=8'h81;
        mem_25[128]=8'h9b;
        mem_25[129]=8'h98;
        mem_25[130]=8'h9d;
        mem_25[131]=8'h9e;
        mem_25[132]=8'h97;
        mem_25[133]=8'h94;
        mem_25[134]=8'h91;
        mem_25[135]=8'h92;
        mem_25[136]=8'h83;
        mem_25[137]=8'h80;
        mem_25[138]=8'h85;
        mem_25[139]=8'h86;
        mem_25[140]=8'h8f;
        mem_25[141]=8'h8c;
        mem_25[142]=8'h89;
        mem_25[143]=8'h8a;
        mem_25[144]=8'hab;
        mem_25[145]=8'ha8;
        mem_25[146]=8'had;
        mem_25[147]=8'hae;
        mem_25[148]=8'ha7;
        mem_25[149]=8'ha4;
        mem_25[150]=8'ha1;
        mem_25[151]=8'ha2;
        mem_25[152]=8'hb3;
        mem_25[153]=8'hb0;
        mem_25[154]=8'hb5;
        mem_25[155]=8'hb6;
        mem_25[156]=8'hbf;
        mem_25[157]=8'hbc;
        mem_25[158]=8'hb9;
        mem_25[159]=8'hba;
        mem_25[160]=8'hfb;
        mem_25[161]=8'hf8;
        mem_25[162]=8'hfd;
        mem_25[163]=8'hfe;
        mem_25[164]=8'hf7;
        mem_25[165]=8'hf4;
        mem_25[166]=8'hf1;
        mem_25[167]=8'hf2;
        mem_25[168]=8'he3;
        mem_25[169]=8'he0;
        mem_25[170]=8'he5;
        mem_25[171]=8'he6;
        mem_25[172]=8'hef;
        mem_25[173]=8'hec;
        mem_25[174]=8'he9;
        mem_25[175]=8'hea;
        mem_25[176]=8'hcb;
        mem_25[177]=8'hc8;
        mem_25[178]=8'hcd;
        mem_25[179]=8'hce;
        mem_25[180]=8'hc7;
        mem_25[181]=8'hc4;
        mem_25[182]=8'hc1;
        mem_25[183]=8'hc2;
        mem_25[184]=8'hd3;
        mem_25[185]=8'hd0;
        mem_25[186]=8'hd5;
        mem_25[187]=8'hd6;
        mem_25[188]=8'hdf;
        mem_25[189]=8'hdc;
        mem_25[190]=8'hd9;
        mem_25[191]=8'hda;
        mem_25[192]=8'h5b;
        mem_25[193]=8'h58;
        mem_25[194]=8'h5d;
        mem_25[195]=8'h5e;
        mem_25[196]=8'h57;
        mem_25[197]=8'h54;
        mem_25[198]=8'h51;
        mem_25[199]=8'h52;
        mem_25[200]=8'h43;
        mem_25[201]=8'h40;
        mem_25[202]=8'h45;
        mem_25[203]=8'h46;
        mem_25[204]=8'h4f;
        mem_25[205]=8'h4c;
        mem_25[206]=8'h49;
        mem_25[207]=8'h4a;
        mem_25[208]=8'h6b;
        mem_25[209]=8'h68;
        mem_25[210]=8'h6d;
        mem_25[211]=8'h6e;
        mem_25[212]=8'h67;
        mem_25[213]=8'h64;
        mem_25[214]=8'h61;
        mem_25[215]=8'h62;
        mem_25[216]=8'h73;
        mem_25[217]=8'h70;
        mem_25[218]=8'h75;
        mem_25[219]=8'h76;
        mem_25[220]=8'h7f;
        mem_25[221]=8'h7c;
        mem_25[222]=8'h79;
        mem_25[223]=8'h7a;
        mem_25[224]=8'h3b;
        mem_25[225]=8'h38;
        mem_25[226]=8'h3d;
        mem_25[227]=8'h3e;
        mem_25[228]=8'h37;
        mem_25[229]=8'h34;
        mem_25[230]=8'h31;
        mem_25[231]=8'h32;
        mem_25[232]=8'h23;
        mem_25[233]=8'h20;
        mem_25[234]=8'h25;
        mem_25[235]=8'h26;
        mem_25[236]=8'h2f;
        mem_25[237]=8'h2c;
        mem_25[238]=8'h29;
        mem_25[239]=8'h2a;
        mem_25[240]=8'hb;
        mem_25[241]=8'h8;
        mem_25[242]=8'hd;
        mem_25[243]=8'he;
        mem_25[244]=8'h7;
        mem_25[245]=8'h4;
        mem_25[246]=8'h1;
        mem_25[247]=8'h2;
        mem_25[248]=8'h13;
        mem_25[249]=8'h10;
        mem_25[250]=8'h15;
        mem_25[251]=8'h16;
        mem_25[252]=8'h1f;
        mem_25[253]=8'h1c;
        mem_25[254]=8'h19;
        mem_25[255]=8'h1a;
    end

    initial begin
        mem_26[0]=8'h0;
        mem_26[1]=8'h2;
        mem_26[2]=8'h4;
        mem_26[3]=8'h6;
        mem_26[4]=8'h8;
        mem_26[5]=8'ha;
        mem_26[6]=8'hc;
        mem_26[7]=8'he;
        mem_26[8]=8'h10;
        mem_26[9]=8'h12;
        mem_26[10]=8'h14;
        mem_26[11]=8'h16;
        mem_26[12]=8'h18;
        mem_26[13]=8'h1a;
        mem_26[14]=8'h1c;
        mem_26[15]=8'h1e;
        mem_26[16]=8'h20;
        mem_26[17]=8'h22;
        mem_26[18]=8'h24;
        mem_26[19]=8'h26;
        mem_26[20]=8'h28;
        mem_26[21]=8'h2a;
        mem_26[22]=8'h2c;
        mem_26[23]=8'h2e;
        mem_26[24]=8'h30;
        mem_26[25]=8'h32;
        mem_26[26]=8'h34;
        mem_26[27]=8'h36;
        mem_26[28]=8'h38;
        mem_26[29]=8'h3a;
        mem_26[30]=8'h3c;
        mem_26[31]=8'h3e;
        mem_26[32]=8'h40;
        mem_26[33]=8'h42;
        mem_26[34]=8'h44;
        mem_26[35]=8'h46;
        mem_26[36]=8'h48;
        mem_26[37]=8'h4a;
        mem_26[38]=8'h4c;
        mem_26[39]=8'h4e;
        mem_26[40]=8'h50;
        mem_26[41]=8'h52;
        mem_26[42]=8'h54;
        mem_26[43]=8'h56;
        mem_26[44]=8'h58;
        mem_26[45]=8'h5a;
        mem_26[46]=8'h5c;
        mem_26[47]=8'h5e;
        mem_26[48]=8'h60;
        mem_26[49]=8'h62;
        mem_26[50]=8'h64;
        mem_26[51]=8'h66;
        mem_26[52]=8'h68;
        mem_26[53]=8'h6a;
        mem_26[54]=8'h6c;
        mem_26[55]=8'h6e;
        mem_26[56]=8'h70;
        mem_26[57]=8'h72;
        mem_26[58]=8'h74;
        mem_26[59]=8'h76;
        mem_26[60]=8'h78;
        mem_26[61]=8'h7a;
        mem_26[62]=8'h7c;
        mem_26[63]=8'h7e;
        mem_26[64]=8'h80;
        mem_26[65]=8'h82;
        mem_26[66]=8'h84;
        mem_26[67]=8'h86;
        mem_26[68]=8'h88;
        mem_26[69]=8'h8a;
        mem_26[70]=8'h8c;
        mem_26[71]=8'h8e;
        mem_26[72]=8'h90;
        mem_26[73]=8'h92;
        mem_26[74]=8'h94;
        mem_26[75]=8'h96;
        mem_26[76]=8'h98;
        mem_26[77]=8'h9a;
        mem_26[78]=8'h9c;
        mem_26[79]=8'h9e;
        mem_26[80]=8'ha0;
        mem_26[81]=8'ha2;
        mem_26[82]=8'ha4;
        mem_26[83]=8'ha6;
        mem_26[84]=8'ha8;
        mem_26[85]=8'haa;
        mem_26[86]=8'hac;
        mem_26[87]=8'hae;
        mem_26[88]=8'hb0;
        mem_26[89]=8'hb2;
        mem_26[90]=8'hb4;
        mem_26[91]=8'hb6;
        mem_26[92]=8'hb8;
        mem_26[93]=8'hba;
        mem_26[94]=8'hbc;
        mem_26[95]=8'hbe;
        mem_26[96]=8'hc0;
        mem_26[97]=8'hc2;
        mem_26[98]=8'hc4;
        mem_26[99]=8'hc6;
        mem_26[100]=8'hc8;
        mem_26[101]=8'hca;
        mem_26[102]=8'hcc;
        mem_26[103]=8'hce;
        mem_26[104]=8'hd0;
        mem_26[105]=8'hd2;
        mem_26[106]=8'hd4;
        mem_26[107]=8'hd6;
        mem_26[108]=8'hd8;
        mem_26[109]=8'hda;
        mem_26[110]=8'hdc;
        mem_26[111]=8'hde;
        mem_26[112]=8'he0;
        mem_26[113]=8'he2;
        mem_26[114]=8'he4;
        mem_26[115]=8'he6;
        mem_26[116]=8'he8;
        mem_26[117]=8'hea;
        mem_26[118]=8'hec;
        mem_26[119]=8'hee;
        mem_26[120]=8'hf0;
        mem_26[121]=8'hf2;
        mem_26[122]=8'hf4;
        mem_26[123]=8'hf6;
        mem_26[124]=8'hf8;
        mem_26[125]=8'hfa;
        mem_26[126]=8'hfc;
        mem_26[127]=8'hfe;
        mem_26[128]=8'h1b;
        mem_26[129]=8'h19;
        mem_26[130]=8'h1f;
        mem_26[131]=8'h1d;
        mem_26[132]=8'h13;
        mem_26[133]=8'h11;
        mem_26[134]=8'h17;
        mem_26[135]=8'h15;
        mem_26[136]=8'hb;
        mem_26[137]=8'h9;
        mem_26[138]=8'hf;
        mem_26[139]=8'hd;
        mem_26[140]=8'h3;
        mem_26[141]=8'h1;
        mem_26[142]=8'h7;
        mem_26[143]=8'h5;
        mem_26[144]=8'h3b;
        mem_26[145]=8'h39;
        mem_26[146]=8'h3f;
        mem_26[147]=8'h3d;
        mem_26[148]=8'h33;
        mem_26[149]=8'h31;
        mem_26[150]=8'h37;
        mem_26[151]=8'h35;
        mem_26[152]=8'h2b;
        mem_26[153]=8'h29;
        mem_26[154]=8'h2f;
        mem_26[155]=8'h2d;
        mem_26[156]=8'h23;
        mem_26[157]=8'h21;
        mem_26[158]=8'h27;
        mem_26[159]=8'h25;
        mem_26[160]=8'h5b;
        mem_26[161]=8'h59;
        mem_26[162]=8'h5f;
        mem_26[163]=8'h5d;
        mem_26[164]=8'h53;
        mem_26[165]=8'h51;
        mem_26[166]=8'h57;
        mem_26[167]=8'h55;
        mem_26[168]=8'h4b;
        mem_26[169]=8'h49;
        mem_26[170]=8'h4f;
        mem_26[171]=8'h4d;
        mem_26[172]=8'h43;
        mem_26[173]=8'h41;
        mem_26[174]=8'h47;
        mem_26[175]=8'h45;
        mem_26[176]=8'h7b;
        mem_26[177]=8'h79;
        mem_26[178]=8'h7f;
        mem_26[179]=8'h7d;
        mem_26[180]=8'h73;
        mem_26[181]=8'h71;
        mem_26[182]=8'h77;
        mem_26[183]=8'h75;
        mem_26[184]=8'h6b;
        mem_26[185]=8'h69;
        mem_26[186]=8'h6f;
        mem_26[187]=8'h6d;
        mem_26[188]=8'h63;
        mem_26[189]=8'h61;
        mem_26[190]=8'h67;
        mem_26[191]=8'h65;
        mem_26[192]=8'h9b;
        mem_26[193]=8'h99;
        mem_26[194]=8'h9f;
        mem_26[195]=8'h9d;
        mem_26[196]=8'h93;
        mem_26[197]=8'h91;
        mem_26[198]=8'h97;
        mem_26[199]=8'h95;
        mem_26[200]=8'h8b;
        mem_26[201]=8'h89;
        mem_26[202]=8'h8f;
        mem_26[203]=8'h8d;
        mem_26[204]=8'h83;
        mem_26[205]=8'h81;
        mem_26[206]=8'h87;
        mem_26[207]=8'h85;
        mem_26[208]=8'hbb;
        mem_26[209]=8'hb9;
        mem_26[210]=8'hbf;
        mem_26[211]=8'hbd;
        mem_26[212]=8'hb3;
        mem_26[213]=8'hb1;
        mem_26[214]=8'hb7;
        mem_26[215]=8'hb5;
        mem_26[216]=8'hab;
        mem_26[217]=8'ha9;
        mem_26[218]=8'haf;
        mem_26[219]=8'had;
        mem_26[220]=8'ha3;
        mem_26[221]=8'ha1;
        mem_26[222]=8'ha7;
        mem_26[223]=8'ha5;
        mem_26[224]=8'hdb;
        mem_26[225]=8'hd9;
        mem_26[226]=8'hdf;
        mem_26[227]=8'hdd;
        mem_26[228]=8'hd3;
        mem_26[229]=8'hd1;
        mem_26[230]=8'hd7;
        mem_26[231]=8'hd5;
        mem_26[232]=8'hcb;
        mem_26[233]=8'hc9;
        mem_26[234]=8'hcf;
        mem_26[235]=8'hcd;
        mem_26[236]=8'hc3;
        mem_26[237]=8'hc1;
        mem_26[238]=8'hc7;
        mem_26[239]=8'hc5;
        mem_26[240]=8'hfb;
        mem_26[241]=8'hf9;
        mem_26[242]=8'hff;
        mem_26[243]=8'hfd;
        mem_26[244]=8'hf3;
        mem_26[245]=8'hf1;
        mem_26[246]=8'hf7;
        mem_26[247]=8'hf5;
        mem_26[248]=8'heb;
        mem_26[249]=8'he9;
        mem_26[250]=8'hef;
        mem_26[251]=8'hed;
        mem_26[252]=8'he3;
        mem_26[253]=8'he1;
        mem_26[254]=8'he7;
        mem_26[255]=8'he5;
    end

    initial begin
        mem_27[0]=8'h0;
        mem_27[1]=8'h3;
        mem_27[2]=8'h6;
        mem_27[3]=8'h5;
        mem_27[4]=8'hc;
        mem_27[5]=8'hf;
        mem_27[6]=8'ha;
        mem_27[7]=8'h9;
        mem_27[8]=8'h18;
        mem_27[9]=8'h1b;
        mem_27[10]=8'h1e;
        mem_27[11]=8'h1d;
        mem_27[12]=8'h14;
        mem_27[13]=8'h17;
        mem_27[14]=8'h12;
        mem_27[15]=8'h11;
        mem_27[16]=8'h30;
        mem_27[17]=8'h33;
        mem_27[18]=8'h36;
        mem_27[19]=8'h35;
        mem_27[20]=8'h3c;
        mem_27[21]=8'h3f;
        mem_27[22]=8'h3a;
        mem_27[23]=8'h39;
        mem_27[24]=8'h28;
        mem_27[25]=8'h2b;
        mem_27[26]=8'h2e;
        mem_27[27]=8'h2d;
        mem_27[28]=8'h24;
        mem_27[29]=8'h27;
        mem_27[30]=8'h22;
        mem_27[31]=8'h21;
        mem_27[32]=8'h60;
        mem_27[33]=8'h63;
        mem_27[34]=8'h66;
        mem_27[35]=8'h65;
        mem_27[36]=8'h6c;
        mem_27[37]=8'h6f;
        mem_27[38]=8'h6a;
        mem_27[39]=8'h69;
        mem_27[40]=8'h78;
        mem_27[41]=8'h7b;
        mem_27[42]=8'h7e;
        mem_27[43]=8'h7d;
        mem_27[44]=8'h74;
        mem_27[45]=8'h77;
        mem_27[46]=8'h72;
        mem_27[47]=8'h71;
        mem_27[48]=8'h50;
        mem_27[49]=8'h53;
        mem_27[50]=8'h56;
        mem_27[51]=8'h55;
        mem_27[52]=8'h5c;
        mem_27[53]=8'h5f;
        mem_27[54]=8'h5a;
        mem_27[55]=8'h59;
        mem_27[56]=8'h48;
        mem_27[57]=8'h4b;
        mem_27[58]=8'h4e;
        mem_27[59]=8'h4d;
        mem_27[60]=8'h44;
        mem_27[61]=8'h47;
        mem_27[62]=8'h42;
        mem_27[63]=8'h41;
        mem_27[64]=8'hc0;
        mem_27[65]=8'hc3;
        mem_27[66]=8'hc6;
        mem_27[67]=8'hc5;
        mem_27[68]=8'hcc;
        mem_27[69]=8'hcf;
        mem_27[70]=8'hca;
        mem_27[71]=8'hc9;
        mem_27[72]=8'hd8;
        mem_27[73]=8'hdb;
        mem_27[74]=8'hde;
        mem_27[75]=8'hdd;
        mem_27[76]=8'hd4;
        mem_27[77]=8'hd7;
        mem_27[78]=8'hd2;
        mem_27[79]=8'hd1;
        mem_27[80]=8'hf0;
        mem_27[81]=8'hf3;
        mem_27[82]=8'hf6;
        mem_27[83]=8'hf5;
        mem_27[84]=8'hfc;
        mem_27[85]=8'hff;
        mem_27[86]=8'hfa;
        mem_27[87]=8'hf9;
        mem_27[88]=8'he8;
        mem_27[89]=8'heb;
        mem_27[90]=8'hee;
        mem_27[91]=8'hed;
        mem_27[92]=8'he4;
        mem_27[93]=8'he7;
        mem_27[94]=8'he2;
        mem_27[95]=8'he1;
        mem_27[96]=8'ha0;
        mem_27[97]=8'ha3;
        mem_27[98]=8'ha6;
        mem_27[99]=8'ha5;
        mem_27[100]=8'hac;
        mem_27[101]=8'haf;
        mem_27[102]=8'haa;
        mem_27[103]=8'ha9;
        mem_27[104]=8'hb8;
        mem_27[105]=8'hbb;
        mem_27[106]=8'hbe;
        mem_27[107]=8'hbd;
        mem_27[108]=8'hb4;
        mem_27[109]=8'hb7;
        mem_27[110]=8'hb2;
        mem_27[111]=8'hb1;
        mem_27[112]=8'h90;
        mem_27[113]=8'h93;
        mem_27[114]=8'h96;
        mem_27[115]=8'h95;
        mem_27[116]=8'h9c;
        mem_27[117]=8'h9f;
        mem_27[118]=8'h9a;
        mem_27[119]=8'h99;
        mem_27[120]=8'h88;
        mem_27[121]=8'h8b;
        mem_27[122]=8'h8e;
        mem_27[123]=8'h8d;
        mem_27[124]=8'h84;
        mem_27[125]=8'h87;
        mem_27[126]=8'h82;
        mem_27[127]=8'h81;
        mem_27[128]=8'h9b;
        mem_27[129]=8'h98;
        mem_27[130]=8'h9d;
        mem_27[131]=8'h9e;
        mem_27[132]=8'h97;
        mem_27[133]=8'h94;
        mem_27[134]=8'h91;
        mem_27[135]=8'h92;
        mem_27[136]=8'h83;
        mem_27[137]=8'h80;
        mem_27[138]=8'h85;
        mem_27[139]=8'h86;
        mem_27[140]=8'h8f;
        mem_27[141]=8'h8c;
        mem_27[142]=8'h89;
        mem_27[143]=8'h8a;
        mem_27[144]=8'hab;
        mem_27[145]=8'ha8;
        mem_27[146]=8'had;
        mem_27[147]=8'hae;
        mem_27[148]=8'ha7;
        mem_27[149]=8'ha4;
        mem_27[150]=8'ha1;
        mem_27[151]=8'ha2;
        mem_27[152]=8'hb3;
        mem_27[153]=8'hb0;
        mem_27[154]=8'hb5;
        mem_27[155]=8'hb6;
        mem_27[156]=8'hbf;
        mem_27[157]=8'hbc;
        mem_27[158]=8'hb9;
        mem_27[159]=8'hba;
        mem_27[160]=8'hfb;
        mem_27[161]=8'hf8;
        mem_27[162]=8'hfd;
        mem_27[163]=8'hfe;
        mem_27[164]=8'hf7;
        mem_27[165]=8'hf4;
        mem_27[166]=8'hf1;
        mem_27[167]=8'hf2;
        mem_27[168]=8'he3;
        mem_27[169]=8'he0;
        mem_27[170]=8'he5;
        mem_27[171]=8'he6;
        mem_27[172]=8'hef;
        mem_27[173]=8'hec;
        mem_27[174]=8'he9;
        mem_27[175]=8'hea;
        mem_27[176]=8'hcb;
        mem_27[177]=8'hc8;
        mem_27[178]=8'hcd;
        mem_27[179]=8'hce;
        mem_27[180]=8'hc7;
        mem_27[181]=8'hc4;
        mem_27[182]=8'hc1;
        mem_27[183]=8'hc2;
        mem_27[184]=8'hd3;
        mem_27[185]=8'hd0;
        mem_27[186]=8'hd5;
        mem_27[187]=8'hd6;
        mem_27[188]=8'hdf;
        mem_27[189]=8'hdc;
        mem_27[190]=8'hd9;
        mem_27[191]=8'hda;
        mem_27[192]=8'h5b;
        mem_27[193]=8'h58;
        mem_27[194]=8'h5d;
        mem_27[195]=8'h5e;
        mem_27[196]=8'h57;
        mem_27[197]=8'h54;
        mem_27[198]=8'h51;
        mem_27[199]=8'h52;
        mem_27[200]=8'h43;
        mem_27[201]=8'h40;
        mem_27[202]=8'h45;
        mem_27[203]=8'h46;
        mem_27[204]=8'h4f;
        mem_27[205]=8'h4c;
        mem_27[206]=8'h49;
        mem_27[207]=8'h4a;
        mem_27[208]=8'h6b;
        mem_27[209]=8'h68;
        mem_27[210]=8'h6d;
        mem_27[211]=8'h6e;
        mem_27[212]=8'h67;
        mem_27[213]=8'h64;
        mem_27[214]=8'h61;
        mem_27[215]=8'h62;
        mem_27[216]=8'h73;
        mem_27[217]=8'h70;
        mem_27[218]=8'h75;
        mem_27[219]=8'h76;
        mem_27[220]=8'h7f;
        mem_27[221]=8'h7c;
        mem_27[222]=8'h79;
        mem_27[223]=8'h7a;
        mem_27[224]=8'h3b;
        mem_27[225]=8'h38;
        mem_27[226]=8'h3d;
        mem_27[227]=8'h3e;
        mem_27[228]=8'h37;
        mem_27[229]=8'h34;
        mem_27[230]=8'h31;
        mem_27[231]=8'h32;
        mem_27[232]=8'h23;
        mem_27[233]=8'h20;
        mem_27[234]=8'h25;
        mem_27[235]=8'h26;
        mem_27[236]=8'h2f;
        mem_27[237]=8'h2c;
        mem_27[238]=8'h29;
        mem_27[239]=8'h2a;
        mem_27[240]=8'hb;
        mem_27[241]=8'h8;
        mem_27[242]=8'hd;
        mem_27[243]=8'he;
        mem_27[244]=8'h7;
        mem_27[245]=8'h4;
        mem_27[246]=8'h1;
        mem_27[247]=8'h2;
        mem_27[248]=8'h13;
        mem_27[249]=8'h10;
        mem_27[250]=8'h15;
        mem_27[251]=8'h16;
        mem_27[252]=8'h1f;
        mem_27[253]=8'h1c;
        mem_27[254]=8'h19;
        mem_27[255]=8'h1a;
    end

    initial begin
        mem_28[0]=8'h0;
        mem_28[1]=8'h2;
        mem_28[2]=8'h4;
        mem_28[3]=8'h6;
        mem_28[4]=8'h8;
        mem_28[5]=8'ha;
        mem_28[6]=8'hc;
        mem_28[7]=8'he;
        mem_28[8]=8'h10;
        mem_28[9]=8'h12;
        mem_28[10]=8'h14;
        mem_28[11]=8'h16;
        mem_28[12]=8'h18;
        mem_28[13]=8'h1a;
        mem_28[14]=8'h1c;
        mem_28[15]=8'h1e;
        mem_28[16]=8'h20;
        mem_28[17]=8'h22;
        mem_28[18]=8'h24;
        mem_28[19]=8'h26;
        mem_28[20]=8'h28;
        mem_28[21]=8'h2a;
        mem_28[22]=8'h2c;
        mem_28[23]=8'h2e;
        mem_28[24]=8'h30;
        mem_28[25]=8'h32;
        mem_28[26]=8'h34;
        mem_28[27]=8'h36;
        mem_28[28]=8'h38;
        mem_28[29]=8'h3a;
        mem_28[30]=8'h3c;
        mem_28[31]=8'h3e;
        mem_28[32]=8'h40;
        mem_28[33]=8'h42;
        mem_28[34]=8'h44;
        mem_28[35]=8'h46;
        mem_28[36]=8'h48;
        mem_28[37]=8'h4a;
        mem_28[38]=8'h4c;
        mem_28[39]=8'h4e;
        mem_28[40]=8'h50;
        mem_28[41]=8'h52;
        mem_28[42]=8'h54;
        mem_28[43]=8'h56;
        mem_28[44]=8'h58;
        mem_28[45]=8'h5a;
        mem_28[46]=8'h5c;
        mem_28[47]=8'h5e;
        mem_28[48]=8'h60;
        mem_28[49]=8'h62;
        mem_28[50]=8'h64;
        mem_28[51]=8'h66;
        mem_28[52]=8'h68;
        mem_28[53]=8'h6a;
        mem_28[54]=8'h6c;
        mem_28[55]=8'h6e;
        mem_28[56]=8'h70;
        mem_28[57]=8'h72;
        mem_28[58]=8'h74;
        mem_28[59]=8'h76;
        mem_28[60]=8'h78;
        mem_28[61]=8'h7a;
        mem_28[62]=8'h7c;
        mem_28[63]=8'h7e;
        mem_28[64]=8'h80;
        mem_28[65]=8'h82;
        mem_28[66]=8'h84;
        mem_28[67]=8'h86;
        mem_28[68]=8'h88;
        mem_28[69]=8'h8a;
        mem_28[70]=8'h8c;
        mem_28[71]=8'h8e;
        mem_28[72]=8'h90;
        mem_28[73]=8'h92;
        mem_28[74]=8'h94;
        mem_28[75]=8'h96;
        mem_28[76]=8'h98;
        mem_28[77]=8'h9a;
        mem_28[78]=8'h9c;
        mem_28[79]=8'h9e;
        mem_28[80]=8'ha0;
        mem_28[81]=8'ha2;
        mem_28[82]=8'ha4;
        mem_28[83]=8'ha6;
        mem_28[84]=8'ha8;
        mem_28[85]=8'haa;
        mem_28[86]=8'hac;
        mem_28[87]=8'hae;
        mem_28[88]=8'hb0;
        mem_28[89]=8'hb2;
        mem_28[90]=8'hb4;
        mem_28[91]=8'hb6;
        mem_28[92]=8'hb8;
        mem_28[93]=8'hba;
        mem_28[94]=8'hbc;
        mem_28[95]=8'hbe;
        mem_28[96]=8'hc0;
        mem_28[97]=8'hc2;
        mem_28[98]=8'hc4;
        mem_28[99]=8'hc6;
        mem_28[100]=8'hc8;
        mem_28[101]=8'hca;
        mem_28[102]=8'hcc;
        mem_28[103]=8'hce;
        mem_28[104]=8'hd0;
        mem_28[105]=8'hd2;
        mem_28[106]=8'hd4;
        mem_28[107]=8'hd6;
        mem_28[108]=8'hd8;
        mem_28[109]=8'hda;
        mem_28[110]=8'hdc;
        mem_28[111]=8'hde;
        mem_28[112]=8'he0;
        mem_28[113]=8'he2;
        mem_28[114]=8'he4;
        mem_28[115]=8'he6;
        mem_28[116]=8'he8;
        mem_28[117]=8'hea;
        mem_28[118]=8'hec;
        mem_28[119]=8'hee;
        mem_28[120]=8'hf0;
        mem_28[121]=8'hf2;
        mem_28[122]=8'hf4;
        mem_28[123]=8'hf6;
        mem_28[124]=8'hf8;
        mem_28[125]=8'hfa;
        mem_28[126]=8'hfc;
        mem_28[127]=8'hfe;
        mem_28[128]=8'h1b;
        mem_28[129]=8'h19;
        mem_28[130]=8'h1f;
        mem_28[131]=8'h1d;
        mem_28[132]=8'h13;
        mem_28[133]=8'h11;
        mem_28[134]=8'h17;
        mem_28[135]=8'h15;
        mem_28[136]=8'hb;
        mem_28[137]=8'h9;
        mem_28[138]=8'hf;
        mem_28[139]=8'hd;
        mem_28[140]=8'h3;
        mem_28[141]=8'h1;
        mem_28[142]=8'h7;
        mem_28[143]=8'h5;
        mem_28[144]=8'h3b;
        mem_28[145]=8'h39;
        mem_28[146]=8'h3f;
        mem_28[147]=8'h3d;
        mem_28[148]=8'h33;
        mem_28[149]=8'h31;
        mem_28[150]=8'h37;
        mem_28[151]=8'h35;
        mem_28[152]=8'h2b;
        mem_28[153]=8'h29;
        mem_28[154]=8'h2f;
        mem_28[155]=8'h2d;
        mem_28[156]=8'h23;
        mem_28[157]=8'h21;
        mem_28[158]=8'h27;
        mem_28[159]=8'h25;
        mem_28[160]=8'h5b;
        mem_28[161]=8'h59;
        mem_28[162]=8'h5f;
        mem_28[163]=8'h5d;
        mem_28[164]=8'h53;
        mem_28[165]=8'h51;
        mem_28[166]=8'h57;
        mem_28[167]=8'h55;
        mem_28[168]=8'h4b;
        mem_28[169]=8'h49;
        mem_28[170]=8'h4f;
        mem_28[171]=8'h4d;
        mem_28[172]=8'h43;
        mem_28[173]=8'h41;
        mem_28[174]=8'h47;
        mem_28[175]=8'h45;
        mem_28[176]=8'h7b;
        mem_28[177]=8'h79;
        mem_28[178]=8'h7f;
        mem_28[179]=8'h7d;
        mem_28[180]=8'h73;
        mem_28[181]=8'h71;
        mem_28[182]=8'h77;
        mem_28[183]=8'h75;
        mem_28[184]=8'h6b;
        mem_28[185]=8'h69;
        mem_28[186]=8'h6f;
        mem_28[187]=8'h6d;
        mem_28[188]=8'h63;
        mem_28[189]=8'h61;
        mem_28[190]=8'h67;
        mem_28[191]=8'h65;
        mem_28[192]=8'h9b;
        mem_28[193]=8'h99;
        mem_28[194]=8'h9f;
        mem_28[195]=8'h9d;
        mem_28[196]=8'h93;
        mem_28[197]=8'h91;
        mem_28[198]=8'h97;
        mem_28[199]=8'h95;
        mem_28[200]=8'h8b;
        mem_28[201]=8'h89;
        mem_28[202]=8'h8f;
        mem_28[203]=8'h8d;
        mem_28[204]=8'h83;
        mem_28[205]=8'h81;
        mem_28[206]=8'h87;
        mem_28[207]=8'h85;
        mem_28[208]=8'hbb;
        mem_28[209]=8'hb9;
        mem_28[210]=8'hbf;
        mem_28[211]=8'hbd;
        mem_28[212]=8'hb3;
        mem_28[213]=8'hb1;
        mem_28[214]=8'hb7;
        mem_28[215]=8'hb5;
        mem_28[216]=8'hab;
        mem_28[217]=8'ha9;
        mem_28[218]=8'haf;
        mem_28[219]=8'had;
        mem_28[220]=8'ha3;
        mem_28[221]=8'ha1;
        mem_28[222]=8'ha7;
        mem_28[223]=8'ha5;
        mem_28[224]=8'hdb;
        mem_28[225]=8'hd9;
        mem_28[226]=8'hdf;
        mem_28[227]=8'hdd;
        mem_28[228]=8'hd3;
        mem_28[229]=8'hd1;
        mem_28[230]=8'hd7;
        mem_28[231]=8'hd5;
        mem_28[232]=8'hcb;
        mem_28[233]=8'hc9;
        mem_28[234]=8'hcf;
        mem_28[235]=8'hcd;
        mem_28[236]=8'hc3;
        mem_28[237]=8'hc1;
        mem_28[238]=8'hc7;
        mem_28[239]=8'hc5;
        mem_28[240]=8'hfb;
        mem_28[241]=8'hf9;
        mem_28[242]=8'hff;
        mem_28[243]=8'hfd;
        mem_28[244]=8'hf3;
        mem_28[245]=8'hf1;
        mem_28[246]=8'hf7;
        mem_28[247]=8'hf5;
        mem_28[248]=8'heb;
        mem_28[249]=8'he9;
        mem_28[250]=8'hef;
        mem_28[251]=8'hed;
        mem_28[252]=8'he3;
        mem_28[253]=8'he1;
        mem_28[254]=8'he7;
        mem_28[255]=8'he5;
    end

    initial begin
        mem_29[0]=8'h0;
        mem_29[1]=8'h3;
        mem_29[2]=8'h6;
        mem_29[3]=8'h5;
        mem_29[4]=8'hc;
        mem_29[5]=8'hf;
        mem_29[6]=8'ha;
        mem_29[7]=8'h9;
        mem_29[8]=8'h18;
        mem_29[9]=8'h1b;
        mem_29[10]=8'h1e;
        mem_29[11]=8'h1d;
        mem_29[12]=8'h14;
        mem_29[13]=8'h17;
        mem_29[14]=8'h12;
        mem_29[15]=8'h11;
        mem_29[16]=8'h30;
        mem_29[17]=8'h33;
        mem_29[18]=8'h36;
        mem_29[19]=8'h35;
        mem_29[20]=8'h3c;
        mem_29[21]=8'h3f;
        mem_29[22]=8'h3a;
        mem_29[23]=8'h39;
        mem_29[24]=8'h28;
        mem_29[25]=8'h2b;
        mem_29[26]=8'h2e;
        mem_29[27]=8'h2d;
        mem_29[28]=8'h24;
        mem_29[29]=8'h27;
        mem_29[30]=8'h22;
        mem_29[31]=8'h21;
        mem_29[32]=8'h60;
        mem_29[33]=8'h63;
        mem_29[34]=8'h66;
        mem_29[35]=8'h65;
        mem_29[36]=8'h6c;
        mem_29[37]=8'h6f;
        mem_29[38]=8'h6a;
        mem_29[39]=8'h69;
        mem_29[40]=8'h78;
        mem_29[41]=8'h7b;
        mem_29[42]=8'h7e;
        mem_29[43]=8'h7d;
        mem_29[44]=8'h74;
        mem_29[45]=8'h77;
        mem_29[46]=8'h72;
        mem_29[47]=8'h71;
        mem_29[48]=8'h50;
        mem_29[49]=8'h53;
        mem_29[50]=8'h56;
        mem_29[51]=8'h55;
        mem_29[52]=8'h5c;
        mem_29[53]=8'h5f;
        mem_29[54]=8'h5a;
        mem_29[55]=8'h59;
        mem_29[56]=8'h48;
        mem_29[57]=8'h4b;
        mem_29[58]=8'h4e;
        mem_29[59]=8'h4d;
        mem_29[60]=8'h44;
        mem_29[61]=8'h47;
        mem_29[62]=8'h42;
        mem_29[63]=8'h41;
        mem_29[64]=8'hc0;
        mem_29[65]=8'hc3;
        mem_29[66]=8'hc6;
        mem_29[67]=8'hc5;
        mem_29[68]=8'hcc;
        mem_29[69]=8'hcf;
        mem_29[70]=8'hca;
        mem_29[71]=8'hc9;
        mem_29[72]=8'hd8;
        mem_29[73]=8'hdb;
        mem_29[74]=8'hde;
        mem_29[75]=8'hdd;
        mem_29[76]=8'hd4;
        mem_29[77]=8'hd7;
        mem_29[78]=8'hd2;
        mem_29[79]=8'hd1;
        mem_29[80]=8'hf0;
        mem_29[81]=8'hf3;
        mem_29[82]=8'hf6;
        mem_29[83]=8'hf5;
        mem_29[84]=8'hfc;
        mem_29[85]=8'hff;
        mem_29[86]=8'hfa;
        mem_29[87]=8'hf9;
        mem_29[88]=8'he8;
        mem_29[89]=8'heb;
        mem_29[90]=8'hee;
        mem_29[91]=8'hed;
        mem_29[92]=8'he4;
        mem_29[93]=8'he7;
        mem_29[94]=8'he2;
        mem_29[95]=8'he1;
        mem_29[96]=8'ha0;
        mem_29[97]=8'ha3;
        mem_29[98]=8'ha6;
        mem_29[99]=8'ha5;
        mem_29[100]=8'hac;
        mem_29[101]=8'haf;
        mem_29[102]=8'haa;
        mem_29[103]=8'ha9;
        mem_29[104]=8'hb8;
        mem_29[105]=8'hbb;
        mem_29[106]=8'hbe;
        mem_29[107]=8'hbd;
        mem_29[108]=8'hb4;
        mem_29[109]=8'hb7;
        mem_29[110]=8'hb2;
        mem_29[111]=8'hb1;
        mem_29[112]=8'h90;
        mem_29[113]=8'h93;
        mem_29[114]=8'h96;
        mem_29[115]=8'h95;
        mem_29[116]=8'h9c;
        mem_29[117]=8'h9f;
        mem_29[118]=8'h9a;
        mem_29[119]=8'h99;
        mem_29[120]=8'h88;
        mem_29[121]=8'h8b;
        mem_29[122]=8'h8e;
        mem_29[123]=8'h8d;
        mem_29[124]=8'h84;
        mem_29[125]=8'h87;
        mem_29[126]=8'h82;
        mem_29[127]=8'h81;
        mem_29[128]=8'h9b;
        mem_29[129]=8'h98;
        mem_29[130]=8'h9d;
        mem_29[131]=8'h9e;
        mem_29[132]=8'h97;
        mem_29[133]=8'h94;
        mem_29[134]=8'h91;
        mem_29[135]=8'h92;
        mem_29[136]=8'h83;
        mem_29[137]=8'h80;
        mem_29[138]=8'h85;
        mem_29[139]=8'h86;
        mem_29[140]=8'h8f;
        mem_29[141]=8'h8c;
        mem_29[142]=8'h89;
        mem_29[143]=8'h8a;
        mem_29[144]=8'hab;
        mem_29[145]=8'ha8;
        mem_29[146]=8'had;
        mem_29[147]=8'hae;
        mem_29[148]=8'ha7;
        mem_29[149]=8'ha4;
        mem_29[150]=8'ha1;
        mem_29[151]=8'ha2;
        mem_29[152]=8'hb3;
        mem_29[153]=8'hb0;
        mem_29[154]=8'hb5;
        mem_29[155]=8'hb6;
        mem_29[156]=8'hbf;
        mem_29[157]=8'hbc;
        mem_29[158]=8'hb9;
        mem_29[159]=8'hba;
        mem_29[160]=8'hfb;
        mem_29[161]=8'hf8;
        mem_29[162]=8'hfd;
        mem_29[163]=8'hfe;
        mem_29[164]=8'hf7;
        mem_29[165]=8'hf4;
        mem_29[166]=8'hf1;
        mem_29[167]=8'hf2;
        mem_29[168]=8'he3;
        mem_29[169]=8'he0;
        mem_29[170]=8'he5;
        mem_29[171]=8'he6;
        mem_29[172]=8'hef;
        mem_29[173]=8'hec;
        mem_29[174]=8'he9;
        mem_29[175]=8'hea;
        mem_29[176]=8'hcb;
        mem_29[177]=8'hc8;
        mem_29[178]=8'hcd;
        mem_29[179]=8'hce;
        mem_29[180]=8'hc7;
        mem_29[181]=8'hc4;
        mem_29[182]=8'hc1;
        mem_29[183]=8'hc2;
        mem_29[184]=8'hd3;
        mem_29[185]=8'hd0;
        mem_29[186]=8'hd5;
        mem_29[187]=8'hd6;
        mem_29[188]=8'hdf;
        mem_29[189]=8'hdc;
        mem_29[190]=8'hd9;
        mem_29[191]=8'hda;
        mem_29[192]=8'h5b;
        mem_29[193]=8'h58;
        mem_29[194]=8'h5d;
        mem_29[195]=8'h5e;
        mem_29[196]=8'h57;
        mem_29[197]=8'h54;
        mem_29[198]=8'h51;
        mem_29[199]=8'h52;
        mem_29[200]=8'h43;
        mem_29[201]=8'h40;
        mem_29[202]=8'h45;
        mem_29[203]=8'h46;
        mem_29[204]=8'h4f;
        mem_29[205]=8'h4c;
        mem_29[206]=8'h49;
        mem_29[207]=8'h4a;
        mem_29[208]=8'h6b;
        mem_29[209]=8'h68;
        mem_29[210]=8'h6d;
        mem_29[211]=8'h6e;
        mem_29[212]=8'h67;
        mem_29[213]=8'h64;
        mem_29[214]=8'h61;
        mem_29[215]=8'h62;
        mem_29[216]=8'h73;
        mem_29[217]=8'h70;
        mem_29[218]=8'h75;
        mem_29[219]=8'h76;
        mem_29[220]=8'h7f;
        mem_29[221]=8'h7c;
        mem_29[222]=8'h79;
        mem_29[223]=8'h7a;
        mem_29[224]=8'h3b;
        mem_29[225]=8'h38;
        mem_29[226]=8'h3d;
        mem_29[227]=8'h3e;
        mem_29[228]=8'h37;
        mem_29[229]=8'h34;
        mem_29[230]=8'h31;
        mem_29[231]=8'h32;
        mem_29[232]=8'h23;
        mem_29[233]=8'h20;
        mem_29[234]=8'h25;
        mem_29[235]=8'h26;
        mem_29[236]=8'h2f;
        mem_29[237]=8'h2c;
        mem_29[238]=8'h29;
        mem_29[239]=8'h2a;
        mem_29[240]=8'hb;
        mem_29[241]=8'h8;
        mem_29[242]=8'hd;
        mem_29[243]=8'he;
        mem_29[244]=8'h7;
        mem_29[245]=8'h4;
        mem_29[246]=8'h1;
        mem_29[247]=8'h2;
        mem_29[248]=8'h13;
        mem_29[249]=8'h10;
        mem_29[250]=8'h15;
        mem_29[251]=8'h16;
        mem_29[252]=8'h1f;
        mem_29[253]=8'h1c;
        mem_29[254]=8'h19;
        mem_29[255]=8'h1a;
    end

    initial begin
        mem_30[0]=8'h0;
        mem_30[1]=8'h2;
        mem_30[2]=8'h4;
        mem_30[3]=8'h6;
        mem_30[4]=8'h8;
        mem_30[5]=8'ha;
        mem_30[6]=8'hc;
        mem_30[7]=8'he;
        mem_30[8]=8'h10;
        mem_30[9]=8'h12;
        mem_30[10]=8'h14;
        mem_30[11]=8'h16;
        mem_30[12]=8'h18;
        mem_30[13]=8'h1a;
        mem_30[14]=8'h1c;
        mem_30[15]=8'h1e;
        mem_30[16]=8'h20;
        mem_30[17]=8'h22;
        mem_30[18]=8'h24;
        mem_30[19]=8'h26;
        mem_30[20]=8'h28;
        mem_30[21]=8'h2a;
        mem_30[22]=8'h2c;
        mem_30[23]=8'h2e;
        mem_30[24]=8'h30;
        mem_30[25]=8'h32;
        mem_30[26]=8'h34;
        mem_30[27]=8'h36;
        mem_30[28]=8'h38;
        mem_30[29]=8'h3a;
        mem_30[30]=8'h3c;
        mem_30[31]=8'h3e;
        mem_30[32]=8'h40;
        mem_30[33]=8'h42;
        mem_30[34]=8'h44;
        mem_30[35]=8'h46;
        mem_30[36]=8'h48;
        mem_30[37]=8'h4a;
        mem_30[38]=8'h4c;
        mem_30[39]=8'h4e;
        mem_30[40]=8'h50;
        mem_30[41]=8'h52;
        mem_30[42]=8'h54;
        mem_30[43]=8'h56;
        mem_30[44]=8'h58;
        mem_30[45]=8'h5a;
        mem_30[46]=8'h5c;
        mem_30[47]=8'h5e;
        mem_30[48]=8'h60;
        mem_30[49]=8'h62;
        mem_30[50]=8'h64;
        mem_30[51]=8'h66;
        mem_30[52]=8'h68;
        mem_30[53]=8'h6a;
        mem_30[54]=8'h6c;
        mem_30[55]=8'h6e;
        mem_30[56]=8'h70;
        mem_30[57]=8'h72;
        mem_30[58]=8'h74;
        mem_30[59]=8'h76;
        mem_30[60]=8'h78;
        mem_30[61]=8'h7a;
        mem_30[62]=8'h7c;
        mem_30[63]=8'h7e;
        mem_30[64]=8'h80;
        mem_30[65]=8'h82;
        mem_30[66]=8'h84;
        mem_30[67]=8'h86;
        mem_30[68]=8'h88;
        mem_30[69]=8'h8a;
        mem_30[70]=8'h8c;
        mem_30[71]=8'h8e;
        mem_30[72]=8'h90;
        mem_30[73]=8'h92;
        mem_30[74]=8'h94;
        mem_30[75]=8'h96;
        mem_30[76]=8'h98;
        mem_30[77]=8'h9a;
        mem_30[78]=8'h9c;
        mem_30[79]=8'h9e;
        mem_30[80]=8'ha0;
        mem_30[81]=8'ha2;
        mem_30[82]=8'ha4;
        mem_30[83]=8'ha6;
        mem_30[84]=8'ha8;
        mem_30[85]=8'haa;
        mem_30[86]=8'hac;
        mem_30[87]=8'hae;
        mem_30[88]=8'hb0;
        mem_30[89]=8'hb2;
        mem_30[90]=8'hb4;
        mem_30[91]=8'hb6;
        mem_30[92]=8'hb8;
        mem_30[93]=8'hba;
        mem_30[94]=8'hbc;
        mem_30[95]=8'hbe;
        mem_30[96]=8'hc0;
        mem_30[97]=8'hc2;
        mem_30[98]=8'hc4;
        mem_30[99]=8'hc6;
        mem_30[100]=8'hc8;
        mem_30[101]=8'hca;
        mem_30[102]=8'hcc;
        mem_30[103]=8'hce;
        mem_30[104]=8'hd0;
        mem_30[105]=8'hd2;
        mem_30[106]=8'hd4;
        mem_30[107]=8'hd6;
        mem_30[108]=8'hd8;
        mem_30[109]=8'hda;
        mem_30[110]=8'hdc;
        mem_30[111]=8'hde;
        mem_30[112]=8'he0;
        mem_30[113]=8'he2;
        mem_30[114]=8'he4;
        mem_30[115]=8'he6;
        mem_30[116]=8'he8;
        mem_30[117]=8'hea;
        mem_30[118]=8'hec;
        mem_30[119]=8'hee;
        mem_30[120]=8'hf0;
        mem_30[121]=8'hf2;
        mem_30[122]=8'hf4;
        mem_30[123]=8'hf6;
        mem_30[124]=8'hf8;
        mem_30[125]=8'hfa;
        mem_30[126]=8'hfc;
        mem_30[127]=8'hfe;
        mem_30[128]=8'h1b;
        mem_30[129]=8'h19;
        mem_30[130]=8'h1f;
        mem_30[131]=8'h1d;
        mem_30[132]=8'h13;
        mem_30[133]=8'h11;
        mem_30[134]=8'h17;
        mem_30[135]=8'h15;
        mem_30[136]=8'hb;
        mem_30[137]=8'h9;
        mem_30[138]=8'hf;
        mem_30[139]=8'hd;
        mem_30[140]=8'h3;
        mem_30[141]=8'h1;
        mem_30[142]=8'h7;
        mem_30[143]=8'h5;
        mem_30[144]=8'h3b;
        mem_30[145]=8'h39;
        mem_30[146]=8'h3f;
        mem_30[147]=8'h3d;
        mem_30[148]=8'h33;
        mem_30[149]=8'h31;
        mem_30[150]=8'h37;
        mem_30[151]=8'h35;
        mem_30[152]=8'h2b;
        mem_30[153]=8'h29;
        mem_30[154]=8'h2f;
        mem_30[155]=8'h2d;
        mem_30[156]=8'h23;
        mem_30[157]=8'h21;
        mem_30[158]=8'h27;
        mem_30[159]=8'h25;
        mem_30[160]=8'h5b;
        mem_30[161]=8'h59;
        mem_30[162]=8'h5f;
        mem_30[163]=8'h5d;
        mem_30[164]=8'h53;
        mem_30[165]=8'h51;
        mem_30[166]=8'h57;
        mem_30[167]=8'h55;
        mem_30[168]=8'h4b;
        mem_30[169]=8'h49;
        mem_30[170]=8'h4f;
        mem_30[171]=8'h4d;
        mem_30[172]=8'h43;
        mem_30[173]=8'h41;
        mem_30[174]=8'h47;
        mem_30[175]=8'h45;
        mem_30[176]=8'h7b;
        mem_30[177]=8'h79;
        mem_30[178]=8'h7f;
        mem_30[179]=8'h7d;
        mem_30[180]=8'h73;
        mem_30[181]=8'h71;
        mem_30[182]=8'h77;
        mem_30[183]=8'h75;
        mem_30[184]=8'h6b;
        mem_30[185]=8'h69;
        mem_30[186]=8'h6f;
        mem_30[187]=8'h6d;
        mem_30[188]=8'h63;
        mem_30[189]=8'h61;
        mem_30[190]=8'h67;
        mem_30[191]=8'h65;
        mem_30[192]=8'h9b;
        mem_30[193]=8'h99;
        mem_30[194]=8'h9f;
        mem_30[195]=8'h9d;
        mem_30[196]=8'h93;
        mem_30[197]=8'h91;
        mem_30[198]=8'h97;
        mem_30[199]=8'h95;
        mem_30[200]=8'h8b;
        mem_30[201]=8'h89;
        mem_30[202]=8'h8f;
        mem_30[203]=8'h8d;
        mem_30[204]=8'h83;
        mem_30[205]=8'h81;
        mem_30[206]=8'h87;
        mem_30[207]=8'h85;
        mem_30[208]=8'hbb;
        mem_30[209]=8'hb9;
        mem_30[210]=8'hbf;
        mem_30[211]=8'hbd;
        mem_30[212]=8'hb3;
        mem_30[213]=8'hb1;
        mem_30[214]=8'hb7;
        mem_30[215]=8'hb5;
        mem_30[216]=8'hab;
        mem_30[217]=8'ha9;
        mem_30[218]=8'haf;
        mem_30[219]=8'had;
        mem_30[220]=8'ha3;
        mem_30[221]=8'ha1;
        mem_30[222]=8'ha7;
        mem_30[223]=8'ha5;
        mem_30[224]=8'hdb;
        mem_30[225]=8'hd9;
        mem_30[226]=8'hdf;
        mem_30[227]=8'hdd;
        mem_30[228]=8'hd3;
        mem_30[229]=8'hd1;
        mem_30[230]=8'hd7;
        mem_30[231]=8'hd5;
        mem_30[232]=8'hcb;
        mem_30[233]=8'hc9;
        mem_30[234]=8'hcf;
        mem_30[235]=8'hcd;
        mem_30[236]=8'hc3;
        mem_30[237]=8'hc1;
        mem_30[238]=8'hc7;
        mem_30[239]=8'hc5;
        mem_30[240]=8'hfb;
        mem_30[241]=8'hf9;
        mem_30[242]=8'hff;
        mem_30[243]=8'hfd;
        mem_30[244]=8'hf3;
        mem_30[245]=8'hf1;
        mem_30[246]=8'hf7;
        mem_30[247]=8'hf5;
        mem_30[248]=8'heb;
        mem_30[249]=8'he9;
        mem_30[250]=8'hef;
        mem_30[251]=8'hed;
        mem_30[252]=8'he3;
        mem_30[253]=8'he1;
        mem_30[254]=8'he7;
        mem_30[255]=8'he5;
    end

    initial begin
        mem_31[0]=8'h0;
        mem_31[1]=8'h3;
        mem_31[2]=8'h6;
        mem_31[3]=8'h5;
        mem_31[4]=8'hc;
        mem_31[5]=8'hf;
        mem_31[6]=8'ha;
        mem_31[7]=8'h9;
        mem_31[8]=8'h18;
        mem_31[9]=8'h1b;
        mem_31[10]=8'h1e;
        mem_31[11]=8'h1d;
        mem_31[12]=8'h14;
        mem_31[13]=8'h17;
        mem_31[14]=8'h12;
        mem_31[15]=8'h11;
        mem_31[16]=8'h30;
        mem_31[17]=8'h33;
        mem_31[18]=8'h36;
        mem_31[19]=8'h35;
        mem_31[20]=8'h3c;
        mem_31[21]=8'h3f;
        mem_31[22]=8'h3a;
        mem_31[23]=8'h39;
        mem_31[24]=8'h28;
        mem_31[25]=8'h2b;
        mem_31[26]=8'h2e;
        mem_31[27]=8'h2d;
        mem_31[28]=8'h24;
        mem_31[29]=8'h27;
        mem_31[30]=8'h22;
        mem_31[31]=8'h21;
        mem_31[32]=8'h60;
        mem_31[33]=8'h63;
        mem_31[34]=8'h66;
        mem_31[35]=8'h65;
        mem_31[36]=8'h6c;
        mem_31[37]=8'h6f;
        mem_31[38]=8'h6a;
        mem_31[39]=8'h69;
        mem_31[40]=8'h78;
        mem_31[41]=8'h7b;
        mem_31[42]=8'h7e;
        mem_31[43]=8'h7d;
        mem_31[44]=8'h74;
        mem_31[45]=8'h77;
        mem_31[46]=8'h72;
        mem_31[47]=8'h71;
        mem_31[48]=8'h50;
        mem_31[49]=8'h53;
        mem_31[50]=8'h56;
        mem_31[51]=8'h55;
        mem_31[52]=8'h5c;
        mem_31[53]=8'h5f;
        mem_31[54]=8'h5a;
        mem_31[55]=8'h59;
        mem_31[56]=8'h48;
        mem_31[57]=8'h4b;
        mem_31[58]=8'h4e;
        mem_31[59]=8'h4d;
        mem_31[60]=8'h44;
        mem_31[61]=8'h47;
        mem_31[62]=8'h42;
        mem_31[63]=8'h41;
        mem_31[64]=8'hc0;
        mem_31[65]=8'hc3;
        mem_31[66]=8'hc6;
        mem_31[67]=8'hc5;
        mem_31[68]=8'hcc;
        mem_31[69]=8'hcf;
        mem_31[70]=8'hca;
        mem_31[71]=8'hc9;
        mem_31[72]=8'hd8;
        mem_31[73]=8'hdb;
        mem_31[74]=8'hde;
        mem_31[75]=8'hdd;
        mem_31[76]=8'hd4;
        mem_31[77]=8'hd7;
        mem_31[78]=8'hd2;
        mem_31[79]=8'hd1;
        mem_31[80]=8'hf0;
        mem_31[81]=8'hf3;
        mem_31[82]=8'hf6;
        mem_31[83]=8'hf5;
        mem_31[84]=8'hfc;
        mem_31[85]=8'hff;
        mem_31[86]=8'hfa;
        mem_31[87]=8'hf9;
        mem_31[88]=8'he8;
        mem_31[89]=8'heb;
        mem_31[90]=8'hee;
        mem_31[91]=8'hed;
        mem_31[92]=8'he4;
        mem_31[93]=8'he7;
        mem_31[94]=8'he2;
        mem_31[95]=8'he1;
        mem_31[96]=8'ha0;
        mem_31[97]=8'ha3;
        mem_31[98]=8'ha6;
        mem_31[99]=8'ha5;
        mem_31[100]=8'hac;
        mem_31[101]=8'haf;
        mem_31[102]=8'haa;
        mem_31[103]=8'ha9;
        mem_31[104]=8'hb8;
        mem_31[105]=8'hbb;
        mem_31[106]=8'hbe;
        mem_31[107]=8'hbd;
        mem_31[108]=8'hb4;
        mem_31[109]=8'hb7;
        mem_31[110]=8'hb2;
        mem_31[111]=8'hb1;
        mem_31[112]=8'h90;
        mem_31[113]=8'h93;
        mem_31[114]=8'h96;
        mem_31[115]=8'h95;
        mem_31[116]=8'h9c;
        mem_31[117]=8'h9f;
        mem_31[118]=8'h9a;
        mem_31[119]=8'h99;
        mem_31[120]=8'h88;
        mem_31[121]=8'h8b;
        mem_31[122]=8'h8e;
        mem_31[123]=8'h8d;
        mem_31[124]=8'h84;
        mem_31[125]=8'h87;
        mem_31[126]=8'h82;
        mem_31[127]=8'h81;
        mem_31[128]=8'h9b;
        mem_31[129]=8'h98;
        mem_31[130]=8'h9d;
        mem_31[131]=8'h9e;
        mem_31[132]=8'h97;
        mem_31[133]=8'h94;
        mem_31[134]=8'h91;
        mem_31[135]=8'h92;
        mem_31[136]=8'h83;
        mem_31[137]=8'h80;
        mem_31[138]=8'h85;
        mem_31[139]=8'h86;
        mem_31[140]=8'h8f;
        mem_31[141]=8'h8c;
        mem_31[142]=8'h89;
        mem_31[143]=8'h8a;
        mem_31[144]=8'hab;
        mem_31[145]=8'ha8;
        mem_31[146]=8'had;
        mem_31[147]=8'hae;
        mem_31[148]=8'ha7;
        mem_31[149]=8'ha4;
        mem_31[150]=8'ha1;
        mem_31[151]=8'ha2;
        mem_31[152]=8'hb3;
        mem_31[153]=8'hb0;
        mem_31[154]=8'hb5;
        mem_31[155]=8'hb6;
        mem_31[156]=8'hbf;
        mem_31[157]=8'hbc;
        mem_31[158]=8'hb9;
        mem_31[159]=8'hba;
        mem_31[160]=8'hfb;
        mem_31[161]=8'hf8;
        mem_31[162]=8'hfd;
        mem_31[163]=8'hfe;
        mem_31[164]=8'hf7;
        mem_31[165]=8'hf4;
        mem_31[166]=8'hf1;
        mem_31[167]=8'hf2;
        mem_31[168]=8'he3;
        mem_31[169]=8'he0;
        mem_31[170]=8'he5;
        mem_31[171]=8'he6;
        mem_31[172]=8'hef;
        mem_31[173]=8'hec;
        mem_31[174]=8'he9;
        mem_31[175]=8'hea;
        mem_31[176]=8'hcb;
        mem_31[177]=8'hc8;
        mem_31[178]=8'hcd;
        mem_31[179]=8'hce;
        mem_31[180]=8'hc7;
        mem_31[181]=8'hc4;
        mem_31[182]=8'hc1;
        mem_31[183]=8'hc2;
        mem_31[184]=8'hd3;
        mem_31[185]=8'hd0;
        mem_31[186]=8'hd5;
        mem_31[187]=8'hd6;
        mem_31[188]=8'hdf;
        mem_31[189]=8'hdc;
        mem_31[190]=8'hd9;
        mem_31[191]=8'hda;
        mem_31[192]=8'h5b;
        mem_31[193]=8'h58;
        mem_31[194]=8'h5d;
        mem_31[195]=8'h5e;
        mem_31[196]=8'h57;
        mem_31[197]=8'h54;
        mem_31[198]=8'h51;
        mem_31[199]=8'h52;
        mem_31[200]=8'h43;
        mem_31[201]=8'h40;
        mem_31[202]=8'h45;
        mem_31[203]=8'h46;
        mem_31[204]=8'h4f;
        mem_31[205]=8'h4c;
        mem_31[206]=8'h49;
        mem_31[207]=8'h4a;
        mem_31[208]=8'h6b;
        mem_31[209]=8'h68;
        mem_31[210]=8'h6d;
        mem_31[211]=8'h6e;
        mem_31[212]=8'h67;
        mem_31[213]=8'h64;
        mem_31[214]=8'h61;
        mem_31[215]=8'h62;
        mem_31[216]=8'h73;
        mem_31[217]=8'h70;
        mem_31[218]=8'h75;
        mem_31[219]=8'h76;
        mem_31[220]=8'h7f;
        mem_31[221]=8'h7c;
        mem_31[222]=8'h79;
        mem_31[223]=8'h7a;
        mem_31[224]=8'h3b;
        mem_31[225]=8'h38;
        mem_31[226]=8'h3d;
        mem_31[227]=8'h3e;
        mem_31[228]=8'h37;
        mem_31[229]=8'h34;
        mem_31[230]=8'h31;
        mem_31[231]=8'h32;
        mem_31[232]=8'h23;
        mem_31[233]=8'h20;
        mem_31[234]=8'h25;
        mem_31[235]=8'h26;
        mem_31[236]=8'h2f;
        mem_31[237]=8'h2c;
        mem_31[238]=8'h29;
        mem_31[239]=8'h2a;
        mem_31[240]=8'hb;
        mem_31[241]=8'h8;
        mem_31[242]=8'hd;
        mem_31[243]=8'he;
        mem_31[244]=8'h7;
        mem_31[245]=8'h4;
        mem_31[246]=8'h1;
        mem_31[247]=8'h2;
        mem_31[248]=8'h13;
        mem_31[249]=8'h10;
        mem_31[250]=8'h15;
        mem_31[251]=8'h16;
        mem_31[252]=8'h1f;
        mem_31[253]=8'h1c;
        mem_31[254]=8'h19;
        mem_31[255]=8'h1a;
    end

    initial begin
        mem_32[0]=8'h0;
        mem_32[1]=8'h2;
        mem_32[2]=8'h4;
        mem_32[3]=8'h6;
        mem_32[4]=8'h8;
        mem_32[5]=8'ha;
        mem_32[6]=8'hc;
        mem_32[7]=8'he;
        mem_32[8]=8'h10;
        mem_32[9]=8'h12;
        mem_32[10]=8'h14;
        mem_32[11]=8'h16;
        mem_32[12]=8'h18;
        mem_32[13]=8'h1a;
        mem_32[14]=8'h1c;
        mem_32[15]=8'h1e;
        mem_32[16]=8'h20;
        mem_32[17]=8'h22;
        mem_32[18]=8'h24;
        mem_32[19]=8'h26;
        mem_32[20]=8'h28;
        mem_32[21]=8'h2a;
        mem_32[22]=8'h2c;
        mem_32[23]=8'h2e;
        mem_32[24]=8'h30;
        mem_32[25]=8'h32;
        mem_32[26]=8'h34;
        mem_32[27]=8'h36;
        mem_32[28]=8'h38;
        mem_32[29]=8'h3a;
        mem_32[30]=8'h3c;
        mem_32[31]=8'h3e;
        mem_32[32]=8'h40;
        mem_32[33]=8'h42;
        mem_32[34]=8'h44;
        mem_32[35]=8'h46;
        mem_32[36]=8'h48;
        mem_32[37]=8'h4a;
        mem_32[38]=8'h4c;
        mem_32[39]=8'h4e;
        mem_32[40]=8'h50;
        mem_32[41]=8'h52;
        mem_32[42]=8'h54;
        mem_32[43]=8'h56;
        mem_32[44]=8'h58;
        mem_32[45]=8'h5a;
        mem_32[46]=8'h5c;
        mem_32[47]=8'h5e;
        mem_32[48]=8'h60;
        mem_32[49]=8'h62;
        mem_32[50]=8'h64;
        mem_32[51]=8'h66;
        mem_32[52]=8'h68;
        mem_32[53]=8'h6a;
        mem_32[54]=8'h6c;
        mem_32[55]=8'h6e;
        mem_32[56]=8'h70;
        mem_32[57]=8'h72;
        mem_32[58]=8'h74;
        mem_32[59]=8'h76;
        mem_32[60]=8'h78;
        mem_32[61]=8'h7a;
        mem_32[62]=8'h7c;
        mem_32[63]=8'h7e;
        mem_32[64]=8'h80;
        mem_32[65]=8'h82;
        mem_32[66]=8'h84;
        mem_32[67]=8'h86;
        mem_32[68]=8'h88;
        mem_32[69]=8'h8a;
        mem_32[70]=8'h8c;
        mem_32[71]=8'h8e;
        mem_32[72]=8'h90;
        mem_32[73]=8'h92;
        mem_32[74]=8'h94;
        mem_32[75]=8'h96;
        mem_32[76]=8'h98;
        mem_32[77]=8'h9a;
        mem_32[78]=8'h9c;
        mem_32[79]=8'h9e;
        mem_32[80]=8'ha0;
        mem_32[81]=8'ha2;
        mem_32[82]=8'ha4;
        mem_32[83]=8'ha6;
        mem_32[84]=8'ha8;
        mem_32[85]=8'haa;
        mem_32[86]=8'hac;
        mem_32[87]=8'hae;
        mem_32[88]=8'hb0;
        mem_32[89]=8'hb2;
        mem_32[90]=8'hb4;
        mem_32[91]=8'hb6;
        mem_32[92]=8'hb8;
        mem_32[93]=8'hba;
        mem_32[94]=8'hbc;
        mem_32[95]=8'hbe;
        mem_32[96]=8'hc0;
        mem_32[97]=8'hc2;
        mem_32[98]=8'hc4;
        mem_32[99]=8'hc6;
        mem_32[100]=8'hc8;
        mem_32[101]=8'hca;
        mem_32[102]=8'hcc;
        mem_32[103]=8'hce;
        mem_32[104]=8'hd0;
        mem_32[105]=8'hd2;
        mem_32[106]=8'hd4;
        mem_32[107]=8'hd6;
        mem_32[108]=8'hd8;
        mem_32[109]=8'hda;
        mem_32[110]=8'hdc;
        mem_32[111]=8'hde;
        mem_32[112]=8'he0;
        mem_32[113]=8'he2;
        mem_32[114]=8'he4;
        mem_32[115]=8'he6;
        mem_32[116]=8'he8;
        mem_32[117]=8'hea;
        mem_32[118]=8'hec;
        mem_32[119]=8'hee;
        mem_32[120]=8'hf0;
        mem_32[121]=8'hf2;
        mem_32[122]=8'hf4;
        mem_32[123]=8'hf6;
        mem_32[124]=8'hf8;
        mem_32[125]=8'hfa;
        mem_32[126]=8'hfc;
        mem_32[127]=8'hfe;
        mem_32[128]=8'h1b;
        mem_32[129]=8'h19;
        mem_32[130]=8'h1f;
        mem_32[131]=8'h1d;
        mem_32[132]=8'h13;
        mem_32[133]=8'h11;
        mem_32[134]=8'h17;
        mem_32[135]=8'h15;
        mem_32[136]=8'hb;
        mem_32[137]=8'h9;
        mem_32[138]=8'hf;
        mem_32[139]=8'hd;
        mem_32[140]=8'h3;
        mem_32[141]=8'h1;
        mem_32[142]=8'h7;
        mem_32[143]=8'h5;
        mem_32[144]=8'h3b;
        mem_32[145]=8'h39;
        mem_32[146]=8'h3f;
        mem_32[147]=8'h3d;
        mem_32[148]=8'h33;
        mem_32[149]=8'h31;
        mem_32[150]=8'h37;
        mem_32[151]=8'h35;
        mem_32[152]=8'h2b;
        mem_32[153]=8'h29;
        mem_32[154]=8'h2f;
        mem_32[155]=8'h2d;
        mem_32[156]=8'h23;
        mem_32[157]=8'h21;
        mem_32[158]=8'h27;
        mem_32[159]=8'h25;
        mem_32[160]=8'h5b;
        mem_32[161]=8'h59;
        mem_32[162]=8'h5f;
        mem_32[163]=8'h5d;
        mem_32[164]=8'h53;
        mem_32[165]=8'h51;
        mem_32[166]=8'h57;
        mem_32[167]=8'h55;
        mem_32[168]=8'h4b;
        mem_32[169]=8'h49;
        mem_32[170]=8'h4f;
        mem_32[171]=8'h4d;
        mem_32[172]=8'h43;
        mem_32[173]=8'h41;
        mem_32[174]=8'h47;
        mem_32[175]=8'h45;
        mem_32[176]=8'h7b;
        mem_32[177]=8'h79;
        mem_32[178]=8'h7f;
        mem_32[179]=8'h7d;
        mem_32[180]=8'h73;
        mem_32[181]=8'h71;
        mem_32[182]=8'h77;
        mem_32[183]=8'h75;
        mem_32[184]=8'h6b;
        mem_32[185]=8'h69;
        mem_32[186]=8'h6f;
        mem_32[187]=8'h6d;
        mem_32[188]=8'h63;
        mem_32[189]=8'h61;
        mem_32[190]=8'h67;
        mem_32[191]=8'h65;
        mem_32[192]=8'h9b;
        mem_32[193]=8'h99;
        mem_32[194]=8'h9f;
        mem_32[195]=8'h9d;
        mem_32[196]=8'h93;
        mem_32[197]=8'h91;
        mem_32[198]=8'h97;
        mem_32[199]=8'h95;
        mem_32[200]=8'h8b;
        mem_32[201]=8'h89;
        mem_32[202]=8'h8f;
        mem_32[203]=8'h8d;
        mem_32[204]=8'h83;
        mem_32[205]=8'h81;
        mem_32[206]=8'h87;
        mem_32[207]=8'h85;
        mem_32[208]=8'hbb;
        mem_32[209]=8'hb9;
        mem_32[210]=8'hbf;
        mem_32[211]=8'hbd;
        mem_32[212]=8'hb3;
        mem_32[213]=8'hb1;
        mem_32[214]=8'hb7;
        mem_32[215]=8'hb5;
        mem_32[216]=8'hab;
        mem_32[217]=8'ha9;
        mem_32[218]=8'haf;
        mem_32[219]=8'had;
        mem_32[220]=8'ha3;
        mem_32[221]=8'ha1;
        mem_32[222]=8'ha7;
        mem_32[223]=8'ha5;
        mem_32[224]=8'hdb;
        mem_32[225]=8'hd9;
        mem_32[226]=8'hdf;
        mem_32[227]=8'hdd;
        mem_32[228]=8'hd3;
        mem_32[229]=8'hd1;
        mem_32[230]=8'hd7;
        mem_32[231]=8'hd5;
        mem_32[232]=8'hcb;
        mem_32[233]=8'hc9;
        mem_32[234]=8'hcf;
        mem_32[235]=8'hcd;
        mem_32[236]=8'hc3;
        mem_32[237]=8'hc1;
        mem_32[238]=8'hc7;
        mem_32[239]=8'hc5;
        mem_32[240]=8'hfb;
        mem_32[241]=8'hf9;
        mem_32[242]=8'hff;
        mem_32[243]=8'hfd;
        mem_32[244]=8'hf3;
        mem_32[245]=8'hf1;
        mem_32[246]=8'hf7;
        mem_32[247]=8'hf5;
        mem_32[248]=8'heb;
        mem_32[249]=8'he9;
        mem_32[250]=8'hef;
        mem_32[251]=8'hed;
        mem_32[252]=8'he3;
        mem_32[253]=8'he1;
        mem_32[254]=8'he7;
        mem_32[255]=8'he5;
    end

    initial begin
        mem_33[0]=8'h0;
        mem_33[1]=8'h3;
        mem_33[2]=8'h6;
        mem_33[3]=8'h5;
        mem_33[4]=8'hc;
        mem_33[5]=8'hf;
        mem_33[6]=8'ha;
        mem_33[7]=8'h9;
        mem_33[8]=8'h18;
        mem_33[9]=8'h1b;
        mem_33[10]=8'h1e;
        mem_33[11]=8'h1d;
        mem_33[12]=8'h14;
        mem_33[13]=8'h17;
        mem_33[14]=8'h12;
        mem_33[15]=8'h11;
        mem_33[16]=8'h30;
        mem_33[17]=8'h33;
        mem_33[18]=8'h36;
        mem_33[19]=8'h35;
        mem_33[20]=8'h3c;
        mem_33[21]=8'h3f;
        mem_33[22]=8'h3a;
        mem_33[23]=8'h39;
        mem_33[24]=8'h28;
        mem_33[25]=8'h2b;
        mem_33[26]=8'h2e;
        mem_33[27]=8'h2d;
        mem_33[28]=8'h24;
        mem_33[29]=8'h27;
        mem_33[30]=8'h22;
        mem_33[31]=8'h21;
        mem_33[32]=8'h60;
        mem_33[33]=8'h63;
        mem_33[34]=8'h66;
        mem_33[35]=8'h65;
        mem_33[36]=8'h6c;
        mem_33[37]=8'h6f;
        mem_33[38]=8'h6a;
        mem_33[39]=8'h69;
        mem_33[40]=8'h78;
        mem_33[41]=8'h7b;
        mem_33[42]=8'h7e;
        mem_33[43]=8'h7d;
        mem_33[44]=8'h74;
        mem_33[45]=8'h77;
        mem_33[46]=8'h72;
        mem_33[47]=8'h71;
        mem_33[48]=8'h50;
        mem_33[49]=8'h53;
        mem_33[50]=8'h56;
        mem_33[51]=8'h55;
        mem_33[52]=8'h5c;
        mem_33[53]=8'h5f;
        mem_33[54]=8'h5a;
        mem_33[55]=8'h59;
        mem_33[56]=8'h48;
        mem_33[57]=8'h4b;
        mem_33[58]=8'h4e;
        mem_33[59]=8'h4d;
        mem_33[60]=8'h44;
        mem_33[61]=8'h47;
        mem_33[62]=8'h42;
        mem_33[63]=8'h41;
        mem_33[64]=8'hc0;
        mem_33[65]=8'hc3;
        mem_33[66]=8'hc6;
        mem_33[67]=8'hc5;
        mem_33[68]=8'hcc;
        mem_33[69]=8'hcf;
        mem_33[70]=8'hca;
        mem_33[71]=8'hc9;
        mem_33[72]=8'hd8;
        mem_33[73]=8'hdb;
        mem_33[74]=8'hde;
        mem_33[75]=8'hdd;
        mem_33[76]=8'hd4;
        mem_33[77]=8'hd7;
        mem_33[78]=8'hd2;
        mem_33[79]=8'hd1;
        mem_33[80]=8'hf0;
        mem_33[81]=8'hf3;
        mem_33[82]=8'hf6;
        mem_33[83]=8'hf5;
        mem_33[84]=8'hfc;
        mem_33[85]=8'hff;
        mem_33[86]=8'hfa;
        mem_33[87]=8'hf9;
        mem_33[88]=8'he8;
        mem_33[89]=8'heb;
        mem_33[90]=8'hee;
        mem_33[91]=8'hed;
        mem_33[92]=8'he4;
        mem_33[93]=8'he7;
        mem_33[94]=8'he2;
        mem_33[95]=8'he1;
        mem_33[96]=8'ha0;
        mem_33[97]=8'ha3;
        mem_33[98]=8'ha6;
        mem_33[99]=8'ha5;
        mem_33[100]=8'hac;
        mem_33[101]=8'haf;
        mem_33[102]=8'haa;
        mem_33[103]=8'ha9;
        mem_33[104]=8'hb8;
        mem_33[105]=8'hbb;
        mem_33[106]=8'hbe;
        mem_33[107]=8'hbd;
        mem_33[108]=8'hb4;
        mem_33[109]=8'hb7;
        mem_33[110]=8'hb2;
        mem_33[111]=8'hb1;
        mem_33[112]=8'h90;
        mem_33[113]=8'h93;
        mem_33[114]=8'h96;
        mem_33[115]=8'h95;
        mem_33[116]=8'h9c;
        mem_33[117]=8'h9f;
        mem_33[118]=8'h9a;
        mem_33[119]=8'h99;
        mem_33[120]=8'h88;
        mem_33[121]=8'h8b;
        mem_33[122]=8'h8e;
        mem_33[123]=8'h8d;
        mem_33[124]=8'h84;
        mem_33[125]=8'h87;
        mem_33[126]=8'h82;
        mem_33[127]=8'h81;
        mem_33[128]=8'h9b;
        mem_33[129]=8'h98;
        mem_33[130]=8'h9d;
        mem_33[131]=8'h9e;
        mem_33[132]=8'h97;
        mem_33[133]=8'h94;
        mem_33[134]=8'h91;
        mem_33[135]=8'h92;
        mem_33[136]=8'h83;
        mem_33[137]=8'h80;
        mem_33[138]=8'h85;
        mem_33[139]=8'h86;
        mem_33[140]=8'h8f;
        mem_33[141]=8'h8c;
        mem_33[142]=8'h89;
        mem_33[143]=8'h8a;
        mem_33[144]=8'hab;
        mem_33[145]=8'ha8;
        mem_33[146]=8'had;
        mem_33[147]=8'hae;
        mem_33[148]=8'ha7;
        mem_33[149]=8'ha4;
        mem_33[150]=8'ha1;
        mem_33[151]=8'ha2;
        mem_33[152]=8'hb3;
        mem_33[153]=8'hb0;
        mem_33[154]=8'hb5;
        mem_33[155]=8'hb6;
        mem_33[156]=8'hbf;
        mem_33[157]=8'hbc;
        mem_33[158]=8'hb9;
        mem_33[159]=8'hba;
        mem_33[160]=8'hfb;
        mem_33[161]=8'hf8;
        mem_33[162]=8'hfd;
        mem_33[163]=8'hfe;
        mem_33[164]=8'hf7;
        mem_33[165]=8'hf4;
        mem_33[166]=8'hf1;
        mem_33[167]=8'hf2;
        mem_33[168]=8'he3;
        mem_33[169]=8'he0;
        mem_33[170]=8'he5;
        mem_33[171]=8'he6;
        mem_33[172]=8'hef;
        mem_33[173]=8'hec;
        mem_33[174]=8'he9;
        mem_33[175]=8'hea;
        mem_33[176]=8'hcb;
        mem_33[177]=8'hc8;
        mem_33[178]=8'hcd;
        mem_33[179]=8'hce;
        mem_33[180]=8'hc7;
        mem_33[181]=8'hc4;
        mem_33[182]=8'hc1;
        mem_33[183]=8'hc2;
        mem_33[184]=8'hd3;
        mem_33[185]=8'hd0;
        mem_33[186]=8'hd5;
        mem_33[187]=8'hd6;
        mem_33[188]=8'hdf;
        mem_33[189]=8'hdc;
        mem_33[190]=8'hd9;
        mem_33[191]=8'hda;
        mem_33[192]=8'h5b;
        mem_33[193]=8'h58;
        mem_33[194]=8'h5d;
        mem_33[195]=8'h5e;
        mem_33[196]=8'h57;
        mem_33[197]=8'h54;
        mem_33[198]=8'h51;
        mem_33[199]=8'h52;
        mem_33[200]=8'h43;
        mem_33[201]=8'h40;
        mem_33[202]=8'h45;
        mem_33[203]=8'h46;
        mem_33[204]=8'h4f;
        mem_33[205]=8'h4c;
        mem_33[206]=8'h49;
        mem_33[207]=8'h4a;
        mem_33[208]=8'h6b;
        mem_33[209]=8'h68;
        mem_33[210]=8'h6d;
        mem_33[211]=8'h6e;
        mem_33[212]=8'h67;
        mem_33[213]=8'h64;
        mem_33[214]=8'h61;
        mem_33[215]=8'h62;
        mem_33[216]=8'h73;
        mem_33[217]=8'h70;
        mem_33[218]=8'h75;
        mem_33[219]=8'h76;
        mem_33[220]=8'h7f;
        mem_33[221]=8'h7c;
        mem_33[222]=8'h79;
        mem_33[223]=8'h7a;
        mem_33[224]=8'h3b;
        mem_33[225]=8'h38;
        mem_33[226]=8'h3d;
        mem_33[227]=8'h3e;
        mem_33[228]=8'h37;
        mem_33[229]=8'h34;
        mem_33[230]=8'h31;
        mem_33[231]=8'h32;
        mem_33[232]=8'h23;
        mem_33[233]=8'h20;
        mem_33[234]=8'h25;
        mem_33[235]=8'h26;
        mem_33[236]=8'h2f;
        mem_33[237]=8'h2c;
        mem_33[238]=8'h29;
        mem_33[239]=8'h2a;
        mem_33[240]=8'hb;
        mem_33[241]=8'h8;
        mem_33[242]=8'hd;
        mem_33[243]=8'he;
        mem_33[244]=8'h7;
        mem_33[245]=8'h4;
        mem_33[246]=8'h1;
        mem_33[247]=8'h2;
        mem_33[248]=8'h13;
        mem_33[249]=8'h10;
        mem_33[250]=8'h15;
        mem_33[251]=8'h16;
        mem_33[252]=8'h1f;
        mem_33[253]=8'h1c;
        mem_33[254]=8'h19;
        mem_33[255]=8'h1a;
    end

    initial begin
        mem_34[0]=8'h0;
        mem_34[1]=8'h2;
        mem_34[2]=8'h4;
        mem_34[3]=8'h6;
        mem_34[4]=8'h8;
        mem_34[5]=8'ha;
        mem_34[6]=8'hc;
        mem_34[7]=8'he;
        mem_34[8]=8'h10;
        mem_34[9]=8'h12;
        mem_34[10]=8'h14;
        mem_34[11]=8'h16;
        mem_34[12]=8'h18;
        mem_34[13]=8'h1a;
        mem_34[14]=8'h1c;
        mem_34[15]=8'h1e;
        mem_34[16]=8'h20;
        mem_34[17]=8'h22;
        mem_34[18]=8'h24;
        mem_34[19]=8'h26;
        mem_34[20]=8'h28;
        mem_34[21]=8'h2a;
        mem_34[22]=8'h2c;
        mem_34[23]=8'h2e;
        mem_34[24]=8'h30;
        mem_34[25]=8'h32;
        mem_34[26]=8'h34;
        mem_34[27]=8'h36;
        mem_34[28]=8'h38;
        mem_34[29]=8'h3a;
        mem_34[30]=8'h3c;
        mem_34[31]=8'h3e;
        mem_34[32]=8'h40;
        mem_34[33]=8'h42;
        mem_34[34]=8'h44;
        mem_34[35]=8'h46;
        mem_34[36]=8'h48;
        mem_34[37]=8'h4a;
        mem_34[38]=8'h4c;
        mem_34[39]=8'h4e;
        mem_34[40]=8'h50;
        mem_34[41]=8'h52;
        mem_34[42]=8'h54;
        mem_34[43]=8'h56;
        mem_34[44]=8'h58;
        mem_34[45]=8'h5a;
        mem_34[46]=8'h5c;
        mem_34[47]=8'h5e;
        mem_34[48]=8'h60;
        mem_34[49]=8'h62;
        mem_34[50]=8'h64;
        mem_34[51]=8'h66;
        mem_34[52]=8'h68;
        mem_34[53]=8'h6a;
        mem_34[54]=8'h6c;
        mem_34[55]=8'h6e;
        mem_34[56]=8'h70;
        mem_34[57]=8'h72;
        mem_34[58]=8'h74;
        mem_34[59]=8'h76;
        mem_34[60]=8'h78;
        mem_34[61]=8'h7a;
        mem_34[62]=8'h7c;
        mem_34[63]=8'h7e;
        mem_34[64]=8'h80;
        mem_34[65]=8'h82;
        mem_34[66]=8'h84;
        mem_34[67]=8'h86;
        mem_34[68]=8'h88;
        mem_34[69]=8'h8a;
        mem_34[70]=8'h8c;
        mem_34[71]=8'h8e;
        mem_34[72]=8'h90;
        mem_34[73]=8'h92;
        mem_34[74]=8'h94;
        mem_34[75]=8'h96;
        mem_34[76]=8'h98;
        mem_34[77]=8'h9a;
        mem_34[78]=8'h9c;
        mem_34[79]=8'h9e;
        mem_34[80]=8'ha0;
        mem_34[81]=8'ha2;
        mem_34[82]=8'ha4;
        mem_34[83]=8'ha6;
        mem_34[84]=8'ha8;
        mem_34[85]=8'haa;
        mem_34[86]=8'hac;
        mem_34[87]=8'hae;
        mem_34[88]=8'hb0;
        mem_34[89]=8'hb2;
        mem_34[90]=8'hb4;
        mem_34[91]=8'hb6;
        mem_34[92]=8'hb8;
        mem_34[93]=8'hba;
        mem_34[94]=8'hbc;
        mem_34[95]=8'hbe;
        mem_34[96]=8'hc0;
        mem_34[97]=8'hc2;
        mem_34[98]=8'hc4;
        mem_34[99]=8'hc6;
        mem_34[100]=8'hc8;
        mem_34[101]=8'hca;
        mem_34[102]=8'hcc;
        mem_34[103]=8'hce;
        mem_34[104]=8'hd0;
        mem_34[105]=8'hd2;
        mem_34[106]=8'hd4;
        mem_34[107]=8'hd6;
        mem_34[108]=8'hd8;
        mem_34[109]=8'hda;
        mem_34[110]=8'hdc;
        mem_34[111]=8'hde;
        mem_34[112]=8'he0;
        mem_34[113]=8'he2;
        mem_34[114]=8'he4;
        mem_34[115]=8'he6;
        mem_34[116]=8'he8;
        mem_34[117]=8'hea;
        mem_34[118]=8'hec;
        mem_34[119]=8'hee;
        mem_34[120]=8'hf0;
        mem_34[121]=8'hf2;
        mem_34[122]=8'hf4;
        mem_34[123]=8'hf6;
        mem_34[124]=8'hf8;
        mem_34[125]=8'hfa;
        mem_34[126]=8'hfc;
        mem_34[127]=8'hfe;
        mem_34[128]=8'h1b;
        mem_34[129]=8'h19;
        mem_34[130]=8'h1f;
        mem_34[131]=8'h1d;
        mem_34[132]=8'h13;
        mem_34[133]=8'h11;
        mem_34[134]=8'h17;
        mem_34[135]=8'h15;
        mem_34[136]=8'hb;
        mem_34[137]=8'h9;
        mem_34[138]=8'hf;
        mem_34[139]=8'hd;
        mem_34[140]=8'h3;
        mem_34[141]=8'h1;
        mem_34[142]=8'h7;
        mem_34[143]=8'h5;
        mem_34[144]=8'h3b;
        mem_34[145]=8'h39;
        mem_34[146]=8'h3f;
        mem_34[147]=8'h3d;
        mem_34[148]=8'h33;
        mem_34[149]=8'h31;
        mem_34[150]=8'h37;
        mem_34[151]=8'h35;
        mem_34[152]=8'h2b;
        mem_34[153]=8'h29;
        mem_34[154]=8'h2f;
        mem_34[155]=8'h2d;
        mem_34[156]=8'h23;
        mem_34[157]=8'h21;
        mem_34[158]=8'h27;
        mem_34[159]=8'h25;
        mem_34[160]=8'h5b;
        mem_34[161]=8'h59;
        mem_34[162]=8'h5f;
        mem_34[163]=8'h5d;
        mem_34[164]=8'h53;
        mem_34[165]=8'h51;
        mem_34[166]=8'h57;
        mem_34[167]=8'h55;
        mem_34[168]=8'h4b;
        mem_34[169]=8'h49;
        mem_34[170]=8'h4f;
        mem_34[171]=8'h4d;
        mem_34[172]=8'h43;
        mem_34[173]=8'h41;
        mem_34[174]=8'h47;
        mem_34[175]=8'h45;
        mem_34[176]=8'h7b;
        mem_34[177]=8'h79;
        mem_34[178]=8'h7f;
        mem_34[179]=8'h7d;
        mem_34[180]=8'h73;
        mem_34[181]=8'h71;
        mem_34[182]=8'h77;
        mem_34[183]=8'h75;
        mem_34[184]=8'h6b;
        mem_34[185]=8'h69;
        mem_34[186]=8'h6f;
        mem_34[187]=8'h6d;
        mem_34[188]=8'h63;
        mem_34[189]=8'h61;
        mem_34[190]=8'h67;
        mem_34[191]=8'h65;
        mem_34[192]=8'h9b;
        mem_34[193]=8'h99;
        mem_34[194]=8'h9f;
        mem_34[195]=8'h9d;
        mem_34[196]=8'h93;
        mem_34[197]=8'h91;
        mem_34[198]=8'h97;
        mem_34[199]=8'h95;
        mem_34[200]=8'h8b;
        mem_34[201]=8'h89;
        mem_34[202]=8'h8f;
        mem_34[203]=8'h8d;
        mem_34[204]=8'h83;
        mem_34[205]=8'h81;
        mem_34[206]=8'h87;
        mem_34[207]=8'h85;
        mem_34[208]=8'hbb;
        mem_34[209]=8'hb9;
        mem_34[210]=8'hbf;
        mem_34[211]=8'hbd;
        mem_34[212]=8'hb3;
        mem_34[213]=8'hb1;
        mem_34[214]=8'hb7;
        mem_34[215]=8'hb5;
        mem_34[216]=8'hab;
        mem_34[217]=8'ha9;
        mem_34[218]=8'haf;
        mem_34[219]=8'had;
        mem_34[220]=8'ha3;
        mem_34[221]=8'ha1;
        mem_34[222]=8'ha7;
        mem_34[223]=8'ha5;
        mem_34[224]=8'hdb;
        mem_34[225]=8'hd9;
        mem_34[226]=8'hdf;
        mem_34[227]=8'hdd;
        mem_34[228]=8'hd3;
        mem_34[229]=8'hd1;
        mem_34[230]=8'hd7;
        mem_34[231]=8'hd5;
        mem_34[232]=8'hcb;
        mem_34[233]=8'hc9;
        mem_34[234]=8'hcf;
        mem_34[235]=8'hcd;
        mem_34[236]=8'hc3;
        mem_34[237]=8'hc1;
        mem_34[238]=8'hc7;
        mem_34[239]=8'hc5;
        mem_34[240]=8'hfb;
        mem_34[241]=8'hf9;
        mem_34[242]=8'hff;
        mem_34[243]=8'hfd;
        mem_34[244]=8'hf3;
        mem_34[245]=8'hf1;
        mem_34[246]=8'hf7;
        mem_34[247]=8'hf5;
        mem_34[248]=8'heb;
        mem_34[249]=8'he9;
        mem_34[250]=8'hef;
        mem_34[251]=8'hed;
        mem_34[252]=8'he3;
        mem_34[253]=8'he1;
        mem_34[254]=8'he7;
        mem_34[255]=8'he5;
    end

    initial begin
        mem_35[0]=8'h0;
        mem_35[1]=8'h3;
        mem_35[2]=8'h6;
        mem_35[3]=8'h5;
        mem_35[4]=8'hc;
        mem_35[5]=8'hf;
        mem_35[6]=8'ha;
        mem_35[7]=8'h9;
        mem_35[8]=8'h18;
        mem_35[9]=8'h1b;
        mem_35[10]=8'h1e;
        mem_35[11]=8'h1d;
        mem_35[12]=8'h14;
        mem_35[13]=8'h17;
        mem_35[14]=8'h12;
        mem_35[15]=8'h11;
        mem_35[16]=8'h30;
        mem_35[17]=8'h33;
        mem_35[18]=8'h36;
        mem_35[19]=8'h35;
        mem_35[20]=8'h3c;
        mem_35[21]=8'h3f;
        mem_35[22]=8'h3a;
        mem_35[23]=8'h39;
        mem_35[24]=8'h28;
        mem_35[25]=8'h2b;
        mem_35[26]=8'h2e;
        mem_35[27]=8'h2d;
        mem_35[28]=8'h24;
        mem_35[29]=8'h27;
        mem_35[30]=8'h22;
        mem_35[31]=8'h21;
        mem_35[32]=8'h60;
        mem_35[33]=8'h63;
        mem_35[34]=8'h66;
        mem_35[35]=8'h65;
        mem_35[36]=8'h6c;
        mem_35[37]=8'h6f;
        mem_35[38]=8'h6a;
        mem_35[39]=8'h69;
        mem_35[40]=8'h78;
        mem_35[41]=8'h7b;
        mem_35[42]=8'h7e;
        mem_35[43]=8'h7d;
        mem_35[44]=8'h74;
        mem_35[45]=8'h77;
        mem_35[46]=8'h72;
        mem_35[47]=8'h71;
        mem_35[48]=8'h50;
        mem_35[49]=8'h53;
        mem_35[50]=8'h56;
        mem_35[51]=8'h55;
        mem_35[52]=8'h5c;
        mem_35[53]=8'h5f;
        mem_35[54]=8'h5a;
        mem_35[55]=8'h59;
        mem_35[56]=8'h48;
        mem_35[57]=8'h4b;
        mem_35[58]=8'h4e;
        mem_35[59]=8'h4d;
        mem_35[60]=8'h44;
        mem_35[61]=8'h47;
        mem_35[62]=8'h42;
        mem_35[63]=8'h41;
        mem_35[64]=8'hc0;
        mem_35[65]=8'hc3;
        mem_35[66]=8'hc6;
        mem_35[67]=8'hc5;
        mem_35[68]=8'hcc;
        mem_35[69]=8'hcf;
        mem_35[70]=8'hca;
        mem_35[71]=8'hc9;
        mem_35[72]=8'hd8;
        mem_35[73]=8'hdb;
        mem_35[74]=8'hde;
        mem_35[75]=8'hdd;
        mem_35[76]=8'hd4;
        mem_35[77]=8'hd7;
        mem_35[78]=8'hd2;
        mem_35[79]=8'hd1;
        mem_35[80]=8'hf0;
        mem_35[81]=8'hf3;
        mem_35[82]=8'hf6;
        mem_35[83]=8'hf5;
        mem_35[84]=8'hfc;
        mem_35[85]=8'hff;
        mem_35[86]=8'hfa;
        mem_35[87]=8'hf9;
        mem_35[88]=8'he8;
        mem_35[89]=8'heb;
        mem_35[90]=8'hee;
        mem_35[91]=8'hed;
        mem_35[92]=8'he4;
        mem_35[93]=8'he7;
        mem_35[94]=8'he2;
        mem_35[95]=8'he1;
        mem_35[96]=8'ha0;
        mem_35[97]=8'ha3;
        mem_35[98]=8'ha6;
        mem_35[99]=8'ha5;
        mem_35[100]=8'hac;
        mem_35[101]=8'haf;
        mem_35[102]=8'haa;
        mem_35[103]=8'ha9;
        mem_35[104]=8'hb8;
        mem_35[105]=8'hbb;
        mem_35[106]=8'hbe;
        mem_35[107]=8'hbd;
        mem_35[108]=8'hb4;
        mem_35[109]=8'hb7;
        mem_35[110]=8'hb2;
        mem_35[111]=8'hb1;
        mem_35[112]=8'h90;
        mem_35[113]=8'h93;
        mem_35[114]=8'h96;
        mem_35[115]=8'h95;
        mem_35[116]=8'h9c;
        mem_35[117]=8'h9f;
        mem_35[118]=8'h9a;
        mem_35[119]=8'h99;
        mem_35[120]=8'h88;
        mem_35[121]=8'h8b;
        mem_35[122]=8'h8e;
        mem_35[123]=8'h8d;
        mem_35[124]=8'h84;
        mem_35[125]=8'h87;
        mem_35[126]=8'h82;
        mem_35[127]=8'h81;
        mem_35[128]=8'h9b;
        mem_35[129]=8'h98;
        mem_35[130]=8'h9d;
        mem_35[131]=8'h9e;
        mem_35[132]=8'h97;
        mem_35[133]=8'h94;
        mem_35[134]=8'h91;
        mem_35[135]=8'h92;
        mem_35[136]=8'h83;
        mem_35[137]=8'h80;
        mem_35[138]=8'h85;
        mem_35[139]=8'h86;
        mem_35[140]=8'h8f;
        mem_35[141]=8'h8c;
        mem_35[142]=8'h89;
        mem_35[143]=8'h8a;
        mem_35[144]=8'hab;
        mem_35[145]=8'ha8;
        mem_35[146]=8'had;
        mem_35[147]=8'hae;
        mem_35[148]=8'ha7;
        mem_35[149]=8'ha4;
        mem_35[150]=8'ha1;
        mem_35[151]=8'ha2;
        mem_35[152]=8'hb3;
        mem_35[153]=8'hb0;
        mem_35[154]=8'hb5;
        mem_35[155]=8'hb6;
        mem_35[156]=8'hbf;
        mem_35[157]=8'hbc;
        mem_35[158]=8'hb9;
        mem_35[159]=8'hba;
        mem_35[160]=8'hfb;
        mem_35[161]=8'hf8;
        mem_35[162]=8'hfd;
        mem_35[163]=8'hfe;
        mem_35[164]=8'hf7;
        mem_35[165]=8'hf4;
        mem_35[166]=8'hf1;
        mem_35[167]=8'hf2;
        mem_35[168]=8'he3;
        mem_35[169]=8'he0;
        mem_35[170]=8'he5;
        mem_35[171]=8'he6;
        mem_35[172]=8'hef;
        mem_35[173]=8'hec;
        mem_35[174]=8'he9;
        mem_35[175]=8'hea;
        mem_35[176]=8'hcb;
        mem_35[177]=8'hc8;
        mem_35[178]=8'hcd;
        mem_35[179]=8'hce;
        mem_35[180]=8'hc7;
        mem_35[181]=8'hc4;
        mem_35[182]=8'hc1;
        mem_35[183]=8'hc2;
        mem_35[184]=8'hd3;
        mem_35[185]=8'hd0;
        mem_35[186]=8'hd5;
        mem_35[187]=8'hd6;
        mem_35[188]=8'hdf;
        mem_35[189]=8'hdc;
        mem_35[190]=8'hd9;
        mem_35[191]=8'hda;
        mem_35[192]=8'h5b;
        mem_35[193]=8'h58;
        mem_35[194]=8'h5d;
        mem_35[195]=8'h5e;
        mem_35[196]=8'h57;
        mem_35[197]=8'h54;
        mem_35[198]=8'h51;
        mem_35[199]=8'h52;
        mem_35[200]=8'h43;
        mem_35[201]=8'h40;
        mem_35[202]=8'h45;
        mem_35[203]=8'h46;
        mem_35[204]=8'h4f;
        mem_35[205]=8'h4c;
        mem_35[206]=8'h49;
        mem_35[207]=8'h4a;
        mem_35[208]=8'h6b;
        mem_35[209]=8'h68;
        mem_35[210]=8'h6d;
        mem_35[211]=8'h6e;
        mem_35[212]=8'h67;
        mem_35[213]=8'h64;
        mem_35[214]=8'h61;
        mem_35[215]=8'h62;
        mem_35[216]=8'h73;
        mem_35[217]=8'h70;
        mem_35[218]=8'h75;
        mem_35[219]=8'h76;
        mem_35[220]=8'h7f;
        mem_35[221]=8'h7c;
        mem_35[222]=8'h79;
        mem_35[223]=8'h7a;
        mem_35[224]=8'h3b;
        mem_35[225]=8'h38;
        mem_35[226]=8'h3d;
        mem_35[227]=8'h3e;
        mem_35[228]=8'h37;
        mem_35[229]=8'h34;
        mem_35[230]=8'h31;
        mem_35[231]=8'h32;
        mem_35[232]=8'h23;
        mem_35[233]=8'h20;
        mem_35[234]=8'h25;
        mem_35[235]=8'h26;
        mem_35[236]=8'h2f;
        mem_35[237]=8'h2c;
        mem_35[238]=8'h29;
        mem_35[239]=8'h2a;
        mem_35[240]=8'hb;
        mem_35[241]=8'h8;
        mem_35[242]=8'hd;
        mem_35[243]=8'he;
        mem_35[244]=8'h7;
        mem_35[245]=8'h4;
        mem_35[246]=8'h1;
        mem_35[247]=8'h2;
        mem_35[248]=8'h13;
        mem_35[249]=8'h10;
        mem_35[250]=8'h15;
        mem_35[251]=8'h16;
        mem_35[252]=8'h1f;
        mem_35[253]=8'h1c;
        mem_35[254]=8'h19;
        mem_35[255]=8'h1a;
    end

    initial begin
        mem_36[0]=8'h0;
        mem_36[1]=8'h2;
        mem_36[2]=8'h4;
        mem_36[3]=8'h6;
        mem_36[4]=8'h8;
        mem_36[5]=8'ha;
        mem_36[6]=8'hc;
        mem_36[7]=8'he;
        mem_36[8]=8'h10;
        mem_36[9]=8'h12;
        mem_36[10]=8'h14;
        mem_36[11]=8'h16;
        mem_36[12]=8'h18;
        mem_36[13]=8'h1a;
        mem_36[14]=8'h1c;
        mem_36[15]=8'h1e;
        mem_36[16]=8'h20;
        mem_36[17]=8'h22;
        mem_36[18]=8'h24;
        mem_36[19]=8'h26;
        mem_36[20]=8'h28;
        mem_36[21]=8'h2a;
        mem_36[22]=8'h2c;
        mem_36[23]=8'h2e;
        mem_36[24]=8'h30;
        mem_36[25]=8'h32;
        mem_36[26]=8'h34;
        mem_36[27]=8'h36;
        mem_36[28]=8'h38;
        mem_36[29]=8'h3a;
        mem_36[30]=8'h3c;
        mem_36[31]=8'h3e;
        mem_36[32]=8'h40;
        mem_36[33]=8'h42;
        mem_36[34]=8'h44;
        mem_36[35]=8'h46;
        mem_36[36]=8'h48;
        mem_36[37]=8'h4a;
        mem_36[38]=8'h4c;
        mem_36[39]=8'h4e;
        mem_36[40]=8'h50;
        mem_36[41]=8'h52;
        mem_36[42]=8'h54;
        mem_36[43]=8'h56;
        mem_36[44]=8'h58;
        mem_36[45]=8'h5a;
        mem_36[46]=8'h5c;
        mem_36[47]=8'h5e;
        mem_36[48]=8'h60;
        mem_36[49]=8'h62;
        mem_36[50]=8'h64;
        mem_36[51]=8'h66;
        mem_36[52]=8'h68;
        mem_36[53]=8'h6a;
        mem_36[54]=8'h6c;
        mem_36[55]=8'h6e;
        mem_36[56]=8'h70;
        mem_36[57]=8'h72;
        mem_36[58]=8'h74;
        mem_36[59]=8'h76;
        mem_36[60]=8'h78;
        mem_36[61]=8'h7a;
        mem_36[62]=8'h7c;
        mem_36[63]=8'h7e;
        mem_36[64]=8'h80;
        mem_36[65]=8'h82;
        mem_36[66]=8'h84;
        mem_36[67]=8'h86;
        mem_36[68]=8'h88;
        mem_36[69]=8'h8a;
        mem_36[70]=8'h8c;
        mem_36[71]=8'h8e;
        mem_36[72]=8'h90;
        mem_36[73]=8'h92;
        mem_36[74]=8'h94;
        mem_36[75]=8'h96;
        mem_36[76]=8'h98;
        mem_36[77]=8'h9a;
        mem_36[78]=8'h9c;
        mem_36[79]=8'h9e;
        mem_36[80]=8'ha0;
        mem_36[81]=8'ha2;
        mem_36[82]=8'ha4;
        mem_36[83]=8'ha6;
        mem_36[84]=8'ha8;
        mem_36[85]=8'haa;
        mem_36[86]=8'hac;
        mem_36[87]=8'hae;
        mem_36[88]=8'hb0;
        mem_36[89]=8'hb2;
        mem_36[90]=8'hb4;
        mem_36[91]=8'hb6;
        mem_36[92]=8'hb8;
        mem_36[93]=8'hba;
        mem_36[94]=8'hbc;
        mem_36[95]=8'hbe;
        mem_36[96]=8'hc0;
        mem_36[97]=8'hc2;
        mem_36[98]=8'hc4;
        mem_36[99]=8'hc6;
        mem_36[100]=8'hc8;
        mem_36[101]=8'hca;
        mem_36[102]=8'hcc;
        mem_36[103]=8'hce;
        mem_36[104]=8'hd0;
        mem_36[105]=8'hd2;
        mem_36[106]=8'hd4;
        mem_36[107]=8'hd6;
        mem_36[108]=8'hd8;
        mem_36[109]=8'hda;
        mem_36[110]=8'hdc;
        mem_36[111]=8'hde;
        mem_36[112]=8'he0;
        mem_36[113]=8'he2;
        mem_36[114]=8'he4;
        mem_36[115]=8'he6;
        mem_36[116]=8'he8;
        mem_36[117]=8'hea;
        mem_36[118]=8'hec;
        mem_36[119]=8'hee;
        mem_36[120]=8'hf0;
        mem_36[121]=8'hf2;
        mem_36[122]=8'hf4;
        mem_36[123]=8'hf6;
        mem_36[124]=8'hf8;
        mem_36[125]=8'hfa;
        mem_36[126]=8'hfc;
        mem_36[127]=8'hfe;
        mem_36[128]=8'h1b;
        mem_36[129]=8'h19;
        mem_36[130]=8'h1f;
        mem_36[131]=8'h1d;
        mem_36[132]=8'h13;
        mem_36[133]=8'h11;
        mem_36[134]=8'h17;
        mem_36[135]=8'h15;
        mem_36[136]=8'hb;
        mem_36[137]=8'h9;
        mem_36[138]=8'hf;
        mem_36[139]=8'hd;
        mem_36[140]=8'h3;
        mem_36[141]=8'h1;
        mem_36[142]=8'h7;
        mem_36[143]=8'h5;
        mem_36[144]=8'h3b;
        mem_36[145]=8'h39;
        mem_36[146]=8'h3f;
        mem_36[147]=8'h3d;
        mem_36[148]=8'h33;
        mem_36[149]=8'h31;
        mem_36[150]=8'h37;
        mem_36[151]=8'h35;
        mem_36[152]=8'h2b;
        mem_36[153]=8'h29;
        mem_36[154]=8'h2f;
        mem_36[155]=8'h2d;
        mem_36[156]=8'h23;
        mem_36[157]=8'h21;
        mem_36[158]=8'h27;
        mem_36[159]=8'h25;
        mem_36[160]=8'h5b;
        mem_36[161]=8'h59;
        mem_36[162]=8'h5f;
        mem_36[163]=8'h5d;
        mem_36[164]=8'h53;
        mem_36[165]=8'h51;
        mem_36[166]=8'h57;
        mem_36[167]=8'h55;
        mem_36[168]=8'h4b;
        mem_36[169]=8'h49;
        mem_36[170]=8'h4f;
        mem_36[171]=8'h4d;
        mem_36[172]=8'h43;
        mem_36[173]=8'h41;
        mem_36[174]=8'h47;
        mem_36[175]=8'h45;
        mem_36[176]=8'h7b;
        mem_36[177]=8'h79;
        mem_36[178]=8'h7f;
        mem_36[179]=8'h7d;
        mem_36[180]=8'h73;
        mem_36[181]=8'h71;
        mem_36[182]=8'h77;
        mem_36[183]=8'h75;
        mem_36[184]=8'h6b;
        mem_36[185]=8'h69;
        mem_36[186]=8'h6f;
        mem_36[187]=8'h6d;
        mem_36[188]=8'h63;
        mem_36[189]=8'h61;
        mem_36[190]=8'h67;
        mem_36[191]=8'h65;
        mem_36[192]=8'h9b;
        mem_36[193]=8'h99;
        mem_36[194]=8'h9f;
        mem_36[195]=8'h9d;
        mem_36[196]=8'h93;
        mem_36[197]=8'h91;
        mem_36[198]=8'h97;
        mem_36[199]=8'h95;
        mem_36[200]=8'h8b;
        mem_36[201]=8'h89;
        mem_36[202]=8'h8f;
        mem_36[203]=8'h8d;
        mem_36[204]=8'h83;
        mem_36[205]=8'h81;
        mem_36[206]=8'h87;
        mem_36[207]=8'h85;
        mem_36[208]=8'hbb;
        mem_36[209]=8'hb9;
        mem_36[210]=8'hbf;
        mem_36[211]=8'hbd;
        mem_36[212]=8'hb3;
        mem_36[213]=8'hb1;
        mem_36[214]=8'hb7;
        mem_36[215]=8'hb5;
        mem_36[216]=8'hab;
        mem_36[217]=8'ha9;
        mem_36[218]=8'haf;
        mem_36[219]=8'had;
        mem_36[220]=8'ha3;
        mem_36[221]=8'ha1;
        mem_36[222]=8'ha7;
        mem_36[223]=8'ha5;
        mem_36[224]=8'hdb;
        mem_36[225]=8'hd9;
        mem_36[226]=8'hdf;
        mem_36[227]=8'hdd;
        mem_36[228]=8'hd3;
        mem_36[229]=8'hd1;
        mem_36[230]=8'hd7;
        mem_36[231]=8'hd5;
        mem_36[232]=8'hcb;
        mem_36[233]=8'hc9;
        mem_36[234]=8'hcf;
        mem_36[235]=8'hcd;
        mem_36[236]=8'hc3;
        mem_36[237]=8'hc1;
        mem_36[238]=8'hc7;
        mem_36[239]=8'hc5;
        mem_36[240]=8'hfb;
        mem_36[241]=8'hf9;
        mem_36[242]=8'hff;
        mem_36[243]=8'hfd;
        mem_36[244]=8'hf3;
        mem_36[245]=8'hf1;
        mem_36[246]=8'hf7;
        mem_36[247]=8'hf5;
        mem_36[248]=8'heb;
        mem_36[249]=8'he9;
        mem_36[250]=8'hef;
        mem_36[251]=8'hed;
        mem_36[252]=8'he3;
        mem_36[253]=8'he1;
        mem_36[254]=8'he7;
        mem_36[255]=8'he5;
    end

    initial begin
        mem_37[0]=8'h0;
        mem_37[1]=8'h3;
        mem_37[2]=8'h6;
        mem_37[3]=8'h5;
        mem_37[4]=8'hc;
        mem_37[5]=8'hf;
        mem_37[6]=8'ha;
        mem_37[7]=8'h9;
        mem_37[8]=8'h18;
        mem_37[9]=8'h1b;
        mem_37[10]=8'h1e;
        mem_37[11]=8'h1d;
        mem_37[12]=8'h14;
        mem_37[13]=8'h17;
        mem_37[14]=8'h12;
        mem_37[15]=8'h11;
        mem_37[16]=8'h30;
        mem_37[17]=8'h33;
        mem_37[18]=8'h36;
        mem_37[19]=8'h35;
        mem_37[20]=8'h3c;
        mem_37[21]=8'h3f;
        mem_37[22]=8'h3a;
        mem_37[23]=8'h39;
        mem_37[24]=8'h28;
        mem_37[25]=8'h2b;
        mem_37[26]=8'h2e;
        mem_37[27]=8'h2d;
        mem_37[28]=8'h24;
        mem_37[29]=8'h27;
        mem_37[30]=8'h22;
        mem_37[31]=8'h21;
        mem_37[32]=8'h60;
        mem_37[33]=8'h63;
        mem_37[34]=8'h66;
        mem_37[35]=8'h65;
        mem_37[36]=8'h6c;
        mem_37[37]=8'h6f;
        mem_37[38]=8'h6a;
        mem_37[39]=8'h69;
        mem_37[40]=8'h78;
        mem_37[41]=8'h7b;
        mem_37[42]=8'h7e;
        mem_37[43]=8'h7d;
        mem_37[44]=8'h74;
        mem_37[45]=8'h77;
        mem_37[46]=8'h72;
        mem_37[47]=8'h71;
        mem_37[48]=8'h50;
        mem_37[49]=8'h53;
        mem_37[50]=8'h56;
        mem_37[51]=8'h55;
        mem_37[52]=8'h5c;
        mem_37[53]=8'h5f;
        mem_37[54]=8'h5a;
        mem_37[55]=8'h59;
        mem_37[56]=8'h48;
        mem_37[57]=8'h4b;
        mem_37[58]=8'h4e;
        mem_37[59]=8'h4d;
        mem_37[60]=8'h44;
        mem_37[61]=8'h47;
        mem_37[62]=8'h42;
        mem_37[63]=8'h41;
        mem_37[64]=8'hc0;
        mem_37[65]=8'hc3;
        mem_37[66]=8'hc6;
        mem_37[67]=8'hc5;
        mem_37[68]=8'hcc;
        mem_37[69]=8'hcf;
        mem_37[70]=8'hca;
        mem_37[71]=8'hc9;
        mem_37[72]=8'hd8;
        mem_37[73]=8'hdb;
        mem_37[74]=8'hde;
        mem_37[75]=8'hdd;
        mem_37[76]=8'hd4;
        mem_37[77]=8'hd7;
        mem_37[78]=8'hd2;
        mem_37[79]=8'hd1;
        mem_37[80]=8'hf0;
        mem_37[81]=8'hf3;
        mem_37[82]=8'hf6;
        mem_37[83]=8'hf5;
        mem_37[84]=8'hfc;
        mem_37[85]=8'hff;
        mem_37[86]=8'hfa;
        mem_37[87]=8'hf9;
        mem_37[88]=8'he8;
        mem_37[89]=8'heb;
        mem_37[90]=8'hee;
        mem_37[91]=8'hed;
        mem_37[92]=8'he4;
        mem_37[93]=8'he7;
        mem_37[94]=8'he2;
        mem_37[95]=8'he1;
        mem_37[96]=8'ha0;
        mem_37[97]=8'ha3;
        mem_37[98]=8'ha6;
        mem_37[99]=8'ha5;
        mem_37[100]=8'hac;
        mem_37[101]=8'haf;
        mem_37[102]=8'haa;
        mem_37[103]=8'ha9;
        mem_37[104]=8'hb8;
        mem_37[105]=8'hbb;
        mem_37[106]=8'hbe;
        mem_37[107]=8'hbd;
        mem_37[108]=8'hb4;
        mem_37[109]=8'hb7;
        mem_37[110]=8'hb2;
        mem_37[111]=8'hb1;
        mem_37[112]=8'h90;
        mem_37[113]=8'h93;
        mem_37[114]=8'h96;
        mem_37[115]=8'h95;
        mem_37[116]=8'h9c;
        mem_37[117]=8'h9f;
        mem_37[118]=8'h9a;
        mem_37[119]=8'h99;
        mem_37[120]=8'h88;
        mem_37[121]=8'h8b;
        mem_37[122]=8'h8e;
        mem_37[123]=8'h8d;
        mem_37[124]=8'h84;
        mem_37[125]=8'h87;
        mem_37[126]=8'h82;
        mem_37[127]=8'h81;
        mem_37[128]=8'h9b;
        mem_37[129]=8'h98;
        mem_37[130]=8'h9d;
        mem_37[131]=8'h9e;
        mem_37[132]=8'h97;
        mem_37[133]=8'h94;
        mem_37[134]=8'h91;
        mem_37[135]=8'h92;
        mem_37[136]=8'h83;
        mem_37[137]=8'h80;
        mem_37[138]=8'h85;
        mem_37[139]=8'h86;
        mem_37[140]=8'h8f;
        mem_37[141]=8'h8c;
        mem_37[142]=8'h89;
        mem_37[143]=8'h8a;
        mem_37[144]=8'hab;
        mem_37[145]=8'ha8;
        mem_37[146]=8'had;
        mem_37[147]=8'hae;
        mem_37[148]=8'ha7;
        mem_37[149]=8'ha4;
        mem_37[150]=8'ha1;
        mem_37[151]=8'ha2;
        mem_37[152]=8'hb3;
        mem_37[153]=8'hb0;
        mem_37[154]=8'hb5;
        mem_37[155]=8'hb6;
        mem_37[156]=8'hbf;
        mem_37[157]=8'hbc;
        mem_37[158]=8'hb9;
        mem_37[159]=8'hba;
        mem_37[160]=8'hfb;
        mem_37[161]=8'hf8;
        mem_37[162]=8'hfd;
        mem_37[163]=8'hfe;
        mem_37[164]=8'hf7;
        mem_37[165]=8'hf4;
        mem_37[166]=8'hf1;
        mem_37[167]=8'hf2;
        mem_37[168]=8'he3;
        mem_37[169]=8'he0;
        mem_37[170]=8'he5;
        mem_37[171]=8'he6;
        mem_37[172]=8'hef;
        mem_37[173]=8'hec;
        mem_37[174]=8'he9;
        mem_37[175]=8'hea;
        mem_37[176]=8'hcb;
        mem_37[177]=8'hc8;
        mem_37[178]=8'hcd;
        mem_37[179]=8'hce;
        mem_37[180]=8'hc7;
        mem_37[181]=8'hc4;
        mem_37[182]=8'hc1;
        mem_37[183]=8'hc2;
        mem_37[184]=8'hd3;
        mem_37[185]=8'hd0;
        mem_37[186]=8'hd5;
        mem_37[187]=8'hd6;
        mem_37[188]=8'hdf;
        mem_37[189]=8'hdc;
        mem_37[190]=8'hd9;
        mem_37[191]=8'hda;
        mem_37[192]=8'h5b;
        mem_37[193]=8'h58;
        mem_37[194]=8'h5d;
        mem_37[195]=8'h5e;
        mem_37[196]=8'h57;
        mem_37[197]=8'h54;
        mem_37[198]=8'h51;
        mem_37[199]=8'h52;
        mem_37[200]=8'h43;
        mem_37[201]=8'h40;
        mem_37[202]=8'h45;
        mem_37[203]=8'h46;
        mem_37[204]=8'h4f;
        mem_37[205]=8'h4c;
        mem_37[206]=8'h49;
        mem_37[207]=8'h4a;
        mem_37[208]=8'h6b;
        mem_37[209]=8'h68;
        mem_37[210]=8'h6d;
        mem_37[211]=8'h6e;
        mem_37[212]=8'h67;
        mem_37[213]=8'h64;
        mem_37[214]=8'h61;
        mem_37[215]=8'h62;
        mem_37[216]=8'h73;
        mem_37[217]=8'h70;
        mem_37[218]=8'h75;
        mem_37[219]=8'h76;
        mem_37[220]=8'h7f;
        mem_37[221]=8'h7c;
        mem_37[222]=8'h79;
        mem_37[223]=8'h7a;
        mem_37[224]=8'h3b;
        mem_37[225]=8'h38;
        mem_37[226]=8'h3d;
        mem_37[227]=8'h3e;
        mem_37[228]=8'h37;
        mem_37[229]=8'h34;
        mem_37[230]=8'h31;
        mem_37[231]=8'h32;
        mem_37[232]=8'h23;
        mem_37[233]=8'h20;
        mem_37[234]=8'h25;
        mem_37[235]=8'h26;
        mem_37[236]=8'h2f;
        mem_37[237]=8'h2c;
        mem_37[238]=8'h29;
        mem_37[239]=8'h2a;
        mem_37[240]=8'hb;
        mem_37[241]=8'h8;
        mem_37[242]=8'hd;
        mem_37[243]=8'he;
        mem_37[244]=8'h7;
        mem_37[245]=8'h4;
        mem_37[246]=8'h1;
        mem_37[247]=8'h2;
        mem_37[248]=8'h13;
        mem_37[249]=8'h10;
        mem_37[250]=8'h15;
        mem_37[251]=8'h16;
        mem_37[252]=8'h1f;
        mem_37[253]=8'h1c;
        mem_37[254]=8'h19;
        mem_37[255]=8'h1a;
    end

    initial begin
        mem_38[0]=8'h0;
        mem_38[1]=8'h2;
        mem_38[2]=8'h4;
        mem_38[3]=8'h6;
        mem_38[4]=8'h8;
        mem_38[5]=8'ha;
        mem_38[6]=8'hc;
        mem_38[7]=8'he;
        mem_38[8]=8'h10;
        mem_38[9]=8'h12;
        mem_38[10]=8'h14;
        mem_38[11]=8'h16;
        mem_38[12]=8'h18;
        mem_38[13]=8'h1a;
        mem_38[14]=8'h1c;
        mem_38[15]=8'h1e;
        mem_38[16]=8'h20;
        mem_38[17]=8'h22;
        mem_38[18]=8'h24;
        mem_38[19]=8'h26;
        mem_38[20]=8'h28;
        mem_38[21]=8'h2a;
        mem_38[22]=8'h2c;
        mem_38[23]=8'h2e;
        mem_38[24]=8'h30;
        mem_38[25]=8'h32;
        mem_38[26]=8'h34;
        mem_38[27]=8'h36;
        mem_38[28]=8'h38;
        mem_38[29]=8'h3a;
        mem_38[30]=8'h3c;
        mem_38[31]=8'h3e;
        mem_38[32]=8'h40;
        mem_38[33]=8'h42;
        mem_38[34]=8'h44;
        mem_38[35]=8'h46;
        mem_38[36]=8'h48;
        mem_38[37]=8'h4a;
        mem_38[38]=8'h4c;
        mem_38[39]=8'h4e;
        mem_38[40]=8'h50;
        mem_38[41]=8'h52;
        mem_38[42]=8'h54;
        mem_38[43]=8'h56;
        mem_38[44]=8'h58;
        mem_38[45]=8'h5a;
        mem_38[46]=8'h5c;
        mem_38[47]=8'h5e;
        mem_38[48]=8'h60;
        mem_38[49]=8'h62;
        mem_38[50]=8'h64;
        mem_38[51]=8'h66;
        mem_38[52]=8'h68;
        mem_38[53]=8'h6a;
        mem_38[54]=8'h6c;
        mem_38[55]=8'h6e;
        mem_38[56]=8'h70;
        mem_38[57]=8'h72;
        mem_38[58]=8'h74;
        mem_38[59]=8'h76;
        mem_38[60]=8'h78;
        mem_38[61]=8'h7a;
        mem_38[62]=8'h7c;
        mem_38[63]=8'h7e;
        mem_38[64]=8'h80;
        mem_38[65]=8'h82;
        mem_38[66]=8'h84;
        mem_38[67]=8'h86;
        mem_38[68]=8'h88;
        mem_38[69]=8'h8a;
        mem_38[70]=8'h8c;
        mem_38[71]=8'h8e;
        mem_38[72]=8'h90;
        mem_38[73]=8'h92;
        mem_38[74]=8'h94;
        mem_38[75]=8'h96;
        mem_38[76]=8'h98;
        mem_38[77]=8'h9a;
        mem_38[78]=8'h9c;
        mem_38[79]=8'h9e;
        mem_38[80]=8'ha0;
        mem_38[81]=8'ha2;
        mem_38[82]=8'ha4;
        mem_38[83]=8'ha6;
        mem_38[84]=8'ha8;
        mem_38[85]=8'haa;
        mem_38[86]=8'hac;
        mem_38[87]=8'hae;
        mem_38[88]=8'hb0;
        mem_38[89]=8'hb2;
        mem_38[90]=8'hb4;
        mem_38[91]=8'hb6;
        mem_38[92]=8'hb8;
        mem_38[93]=8'hba;
        mem_38[94]=8'hbc;
        mem_38[95]=8'hbe;
        mem_38[96]=8'hc0;
        mem_38[97]=8'hc2;
        mem_38[98]=8'hc4;
        mem_38[99]=8'hc6;
        mem_38[100]=8'hc8;
        mem_38[101]=8'hca;
        mem_38[102]=8'hcc;
        mem_38[103]=8'hce;
        mem_38[104]=8'hd0;
        mem_38[105]=8'hd2;
        mem_38[106]=8'hd4;
        mem_38[107]=8'hd6;
        mem_38[108]=8'hd8;
        mem_38[109]=8'hda;
        mem_38[110]=8'hdc;
        mem_38[111]=8'hde;
        mem_38[112]=8'he0;
        mem_38[113]=8'he2;
        mem_38[114]=8'he4;
        mem_38[115]=8'he6;
        mem_38[116]=8'he8;
        mem_38[117]=8'hea;
        mem_38[118]=8'hec;
        mem_38[119]=8'hee;
        mem_38[120]=8'hf0;
        mem_38[121]=8'hf2;
        mem_38[122]=8'hf4;
        mem_38[123]=8'hf6;
        mem_38[124]=8'hf8;
        mem_38[125]=8'hfa;
        mem_38[126]=8'hfc;
        mem_38[127]=8'hfe;
        mem_38[128]=8'h1b;
        mem_38[129]=8'h19;
        mem_38[130]=8'h1f;
        mem_38[131]=8'h1d;
        mem_38[132]=8'h13;
        mem_38[133]=8'h11;
        mem_38[134]=8'h17;
        mem_38[135]=8'h15;
        mem_38[136]=8'hb;
        mem_38[137]=8'h9;
        mem_38[138]=8'hf;
        mem_38[139]=8'hd;
        mem_38[140]=8'h3;
        mem_38[141]=8'h1;
        mem_38[142]=8'h7;
        mem_38[143]=8'h5;
        mem_38[144]=8'h3b;
        mem_38[145]=8'h39;
        mem_38[146]=8'h3f;
        mem_38[147]=8'h3d;
        mem_38[148]=8'h33;
        mem_38[149]=8'h31;
        mem_38[150]=8'h37;
        mem_38[151]=8'h35;
        mem_38[152]=8'h2b;
        mem_38[153]=8'h29;
        mem_38[154]=8'h2f;
        mem_38[155]=8'h2d;
        mem_38[156]=8'h23;
        mem_38[157]=8'h21;
        mem_38[158]=8'h27;
        mem_38[159]=8'h25;
        mem_38[160]=8'h5b;
        mem_38[161]=8'h59;
        mem_38[162]=8'h5f;
        mem_38[163]=8'h5d;
        mem_38[164]=8'h53;
        mem_38[165]=8'h51;
        mem_38[166]=8'h57;
        mem_38[167]=8'h55;
        mem_38[168]=8'h4b;
        mem_38[169]=8'h49;
        mem_38[170]=8'h4f;
        mem_38[171]=8'h4d;
        mem_38[172]=8'h43;
        mem_38[173]=8'h41;
        mem_38[174]=8'h47;
        mem_38[175]=8'h45;
        mem_38[176]=8'h7b;
        mem_38[177]=8'h79;
        mem_38[178]=8'h7f;
        mem_38[179]=8'h7d;
        mem_38[180]=8'h73;
        mem_38[181]=8'h71;
        mem_38[182]=8'h77;
        mem_38[183]=8'h75;
        mem_38[184]=8'h6b;
        mem_38[185]=8'h69;
        mem_38[186]=8'h6f;
        mem_38[187]=8'h6d;
        mem_38[188]=8'h63;
        mem_38[189]=8'h61;
        mem_38[190]=8'h67;
        mem_38[191]=8'h65;
        mem_38[192]=8'h9b;
        mem_38[193]=8'h99;
        mem_38[194]=8'h9f;
        mem_38[195]=8'h9d;
        mem_38[196]=8'h93;
        mem_38[197]=8'h91;
        mem_38[198]=8'h97;
        mem_38[199]=8'h95;
        mem_38[200]=8'h8b;
        mem_38[201]=8'h89;
        mem_38[202]=8'h8f;
        mem_38[203]=8'h8d;
        mem_38[204]=8'h83;
        mem_38[205]=8'h81;
        mem_38[206]=8'h87;
        mem_38[207]=8'h85;
        mem_38[208]=8'hbb;
        mem_38[209]=8'hb9;
        mem_38[210]=8'hbf;
        mem_38[211]=8'hbd;
        mem_38[212]=8'hb3;
        mem_38[213]=8'hb1;
        mem_38[214]=8'hb7;
        mem_38[215]=8'hb5;
        mem_38[216]=8'hab;
        mem_38[217]=8'ha9;
        mem_38[218]=8'haf;
        mem_38[219]=8'had;
        mem_38[220]=8'ha3;
        mem_38[221]=8'ha1;
        mem_38[222]=8'ha7;
        mem_38[223]=8'ha5;
        mem_38[224]=8'hdb;
        mem_38[225]=8'hd9;
        mem_38[226]=8'hdf;
        mem_38[227]=8'hdd;
        mem_38[228]=8'hd3;
        mem_38[229]=8'hd1;
        mem_38[230]=8'hd7;
        mem_38[231]=8'hd5;
        mem_38[232]=8'hcb;
        mem_38[233]=8'hc9;
        mem_38[234]=8'hcf;
        mem_38[235]=8'hcd;
        mem_38[236]=8'hc3;
        mem_38[237]=8'hc1;
        mem_38[238]=8'hc7;
        mem_38[239]=8'hc5;
        mem_38[240]=8'hfb;
        mem_38[241]=8'hf9;
        mem_38[242]=8'hff;
        mem_38[243]=8'hfd;
        mem_38[244]=8'hf3;
        mem_38[245]=8'hf1;
        mem_38[246]=8'hf7;
        mem_38[247]=8'hf5;
        mem_38[248]=8'heb;
        mem_38[249]=8'he9;
        mem_38[250]=8'hef;
        mem_38[251]=8'hed;
        mem_38[252]=8'he3;
        mem_38[253]=8'he1;
        mem_38[254]=8'he7;
        mem_38[255]=8'he5;
    end

    initial begin
        mem_39[0]=8'h0;
        mem_39[1]=8'h3;
        mem_39[2]=8'h6;
        mem_39[3]=8'h5;
        mem_39[4]=8'hc;
        mem_39[5]=8'hf;
        mem_39[6]=8'ha;
        mem_39[7]=8'h9;
        mem_39[8]=8'h18;
        mem_39[9]=8'h1b;
        mem_39[10]=8'h1e;
        mem_39[11]=8'h1d;
        mem_39[12]=8'h14;
        mem_39[13]=8'h17;
        mem_39[14]=8'h12;
        mem_39[15]=8'h11;
        mem_39[16]=8'h30;
        mem_39[17]=8'h33;
        mem_39[18]=8'h36;
        mem_39[19]=8'h35;
        mem_39[20]=8'h3c;
        mem_39[21]=8'h3f;
        mem_39[22]=8'h3a;
        mem_39[23]=8'h39;
        mem_39[24]=8'h28;
        mem_39[25]=8'h2b;
        mem_39[26]=8'h2e;
        mem_39[27]=8'h2d;
        mem_39[28]=8'h24;
        mem_39[29]=8'h27;
        mem_39[30]=8'h22;
        mem_39[31]=8'h21;
        mem_39[32]=8'h60;
        mem_39[33]=8'h63;
        mem_39[34]=8'h66;
        mem_39[35]=8'h65;
        mem_39[36]=8'h6c;
        mem_39[37]=8'h6f;
        mem_39[38]=8'h6a;
        mem_39[39]=8'h69;
        mem_39[40]=8'h78;
        mem_39[41]=8'h7b;
        mem_39[42]=8'h7e;
        mem_39[43]=8'h7d;
        mem_39[44]=8'h74;
        mem_39[45]=8'h77;
        mem_39[46]=8'h72;
        mem_39[47]=8'h71;
        mem_39[48]=8'h50;
        mem_39[49]=8'h53;
        mem_39[50]=8'h56;
        mem_39[51]=8'h55;
        mem_39[52]=8'h5c;
        mem_39[53]=8'h5f;
        mem_39[54]=8'h5a;
        mem_39[55]=8'h59;
        mem_39[56]=8'h48;
        mem_39[57]=8'h4b;
        mem_39[58]=8'h4e;
        mem_39[59]=8'h4d;
        mem_39[60]=8'h44;
        mem_39[61]=8'h47;
        mem_39[62]=8'h42;
        mem_39[63]=8'h41;
        mem_39[64]=8'hc0;
        mem_39[65]=8'hc3;
        mem_39[66]=8'hc6;
        mem_39[67]=8'hc5;
        mem_39[68]=8'hcc;
        mem_39[69]=8'hcf;
        mem_39[70]=8'hca;
        mem_39[71]=8'hc9;
        mem_39[72]=8'hd8;
        mem_39[73]=8'hdb;
        mem_39[74]=8'hde;
        mem_39[75]=8'hdd;
        mem_39[76]=8'hd4;
        mem_39[77]=8'hd7;
        mem_39[78]=8'hd2;
        mem_39[79]=8'hd1;
        mem_39[80]=8'hf0;
        mem_39[81]=8'hf3;
        mem_39[82]=8'hf6;
        mem_39[83]=8'hf5;
        mem_39[84]=8'hfc;
        mem_39[85]=8'hff;
        mem_39[86]=8'hfa;
        mem_39[87]=8'hf9;
        mem_39[88]=8'he8;
        mem_39[89]=8'heb;
        mem_39[90]=8'hee;
        mem_39[91]=8'hed;
        mem_39[92]=8'he4;
        mem_39[93]=8'he7;
        mem_39[94]=8'he2;
        mem_39[95]=8'he1;
        mem_39[96]=8'ha0;
        mem_39[97]=8'ha3;
        mem_39[98]=8'ha6;
        mem_39[99]=8'ha5;
        mem_39[100]=8'hac;
        mem_39[101]=8'haf;
        mem_39[102]=8'haa;
        mem_39[103]=8'ha9;
        mem_39[104]=8'hb8;
        mem_39[105]=8'hbb;
        mem_39[106]=8'hbe;
        mem_39[107]=8'hbd;
        mem_39[108]=8'hb4;
        mem_39[109]=8'hb7;
        mem_39[110]=8'hb2;
        mem_39[111]=8'hb1;
        mem_39[112]=8'h90;
        mem_39[113]=8'h93;
        mem_39[114]=8'h96;
        mem_39[115]=8'h95;
        mem_39[116]=8'h9c;
        mem_39[117]=8'h9f;
        mem_39[118]=8'h9a;
        mem_39[119]=8'h99;
        mem_39[120]=8'h88;
        mem_39[121]=8'h8b;
        mem_39[122]=8'h8e;
        mem_39[123]=8'h8d;
        mem_39[124]=8'h84;
        mem_39[125]=8'h87;
        mem_39[126]=8'h82;
        mem_39[127]=8'h81;
        mem_39[128]=8'h9b;
        mem_39[129]=8'h98;
        mem_39[130]=8'h9d;
        mem_39[131]=8'h9e;
        mem_39[132]=8'h97;
        mem_39[133]=8'h94;
        mem_39[134]=8'h91;
        mem_39[135]=8'h92;
        mem_39[136]=8'h83;
        mem_39[137]=8'h80;
        mem_39[138]=8'h85;
        mem_39[139]=8'h86;
        mem_39[140]=8'h8f;
        mem_39[141]=8'h8c;
        mem_39[142]=8'h89;
        mem_39[143]=8'h8a;
        mem_39[144]=8'hab;
        mem_39[145]=8'ha8;
        mem_39[146]=8'had;
        mem_39[147]=8'hae;
        mem_39[148]=8'ha7;
        mem_39[149]=8'ha4;
        mem_39[150]=8'ha1;
        mem_39[151]=8'ha2;
        mem_39[152]=8'hb3;
        mem_39[153]=8'hb0;
        mem_39[154]=8'hb5;
        mem_39[155]=8'hb6;
        mem_39[156]=8'hbf;
        mem_39[157]=8'hbc;
        mem_39[158]=8'hb9;
        mem_39[159]=8'hba;
        mem_39[160]=8'hfb;
        mem_39[161]=8'hf8;
        mem_39[162]=8'hfd;
        mem_39[163]=8'hfe;
        mem_39[164]=8'hf7;
        mem_39[165]=8'hf4;
        mem_39[166]=8'hf1;
        mem_39[167]=8'hf2;
        mem_39[168]=8'he3;
        mem_39[169]=8'he0;
        mem_39[170]=8'he5;
        mem_39[171]=8'he6;
        mem_39[172]=8'hef;
        mem_39[173]=8'hec;
        mem_39[174]=8'he9;
        mem_39[175]=8'hea;
        mem_39[176]=8'hcb;
        mem_39[177]=8'hc8;
        mem_39[178]=8'hcd;
        mem_39[179]=8'hce;
        mem_39[180]=8'hc7;
        mem_39[181]=8'hc4;
        mem_39[182]=8'hc1;
        mem_39[183]=8'hc2;
        mem_39[184]=8'hd3;
        mem_39[185]=8'hd0;
        mem_39[186]=8'hd5;
        mem_39[187]=8'hd6;
        mem_39[188]=8'hdf;
        mem_39[189]=8'hdc;
        mem_39[190]=8'hd9;
        mem_39[191]=8'hda;
        mem_39[192]=8'h5b;
        mem_39[193]=8'h58;
        mem_39[194]=8'h5d;
        mem_39[195]=8'h5e;
        mem_39[196]=8'h57;
        mem_39[197]=8'h54;
        mem_39[198]=8'h51;
        mem_39[199]=8'h52;
        mem_39[200]=8'h43;
        mem_39[201]=8'h40;
        mem_39[202]=8'h45;
        mem_39[203]=8'h46;
        mem_39[204]=8'h4f;
        mem_39[205]=8'h4c;
        mem_39[206]=8'h49;
        mem_39[207]=8'h4a;
        mem_39[208]=8'h6b;
        mem_39[209]=8'h68;
        mem_39[210]=8'h6d;
        mem_39[211]=8'h6e;
        mem_39[212]=8'h67;
        mem_39[213]=8'h64;
        mem_39[214]=8'h61;
        mem_39[215]=8'h62;
        mem_39[216]=8'h73;
        mem_39[217]=8'h70;
        mem_39[218]=8'h75;
        mem_39[219]=8'h76;
        mem_39[220]=8'h7f;
        mem_39[221]=8'h7c;
        mem_39[222]=8'h79;
        mem_39[223]=8'h7a;
        mem_39[224]=8'h3b;
        mem_39[225]=8'h38;
        mem_39[226]=8'h3d;
        mem_39[227]=8'h3e;
        mem_39[228]=8'h37;
        mem_39[229]=8'h34;
        mem_39[230]=8'h31;
        mem_39[231]=8'h32;
        mem_39[232]=8'h23;
        mem_39[233]=8'h20;
        mem_39[234]=8'h25;
        mem_39[235]=8'h26;
        mem_39[236]=8'h2f;
        mem_39[237]=8'h2c;
        mem_39[238]=8'h29;
        mem_39[239]=8'h2a;
        mem_39[240]=8'hb;
        mem_39[241]=8'h8;
        mem_39[242]=8'hd;
        mem_39[243]=8'he;
        mem_39[244]=8'h7;
        mem_39[245]=8'h4;
        mem_39[246]=8'h1;
        mem_39[247]=8'h2;
        mem_39[248]=8'h13;
        mem_39[249]=8'h10;
        mem_39[250]=8'h15;
        mem_39[251]=8'h16;
        mem_39[252]=8'h1f;
        mem_39[253]=8'h1c;
        mem_39[254]=8'h19;
        mem_39[255]=8'h1a;
    end

    initial begin
        mem_40[0]=8'h0;
        mem_40[1]=8'h2;
        mem_40[2]=8'h4;
        mem_40[3]=8'h6;
        mem_40[4]=8'h8;
        mem_40[5]=8'ha;
        mem_40[6]=8'hc;
        mem_40[7]=8'he;
        mem_40[8]=8'h10;
        mem_40[9]=8'h12;
        mem_40[10]=8'h14;
        mem_40[11]=8'h16;
        mem_40[12]=8'h18;
        mem_40[13]=8'h1a;
        mem_40[14]=8'h1c;
        mem_40[15]=8'h1e;
        mem_40[16]=8'h20;
        mem_40[17]=8'h22;
        mem_40[18]=8'h24;
        mem_40[19]=8'h26;
        mem_40[20]=8'h28;
        mem_40[21]=8'h2a;
        mem_40[22]=8'h2c;
        mem_40[23]=8'h2e;
        mem_40[24]=8'h30;
        mem_40[25]=8'h32;
        mem_40[26]=8'h34;
        mem_40[27]=8'h36;
        mem_40[28]=8'h38;
        mem_40[29]=8'h3a;
        mem_40[30]=8'h3c;
        mem_40[31]=8'h3e;
        mem_40[32]=8'h40;
        mem_40[33]=8'h42;
        mem_40[34]=8'h44;
        mem_40[35]=8'h46;
        mem_40[36]=8'h48;
        mem_40[37]=8'h4a;
        mem_40[38]=8'h4c;
        mem_40[39]=8'h4e;
        mem_40[40]=8'h50;
        mem_40[41]=8'h52;
        mem_40[42]=8'h54;
        mem_40[43]=8'h56;
        mem_40[44]=8'h58;
        mem_40[45]=8'h5a;
        mem_40[46]=8'h5c;
        mem_40[47]=8'h5e;
        mem_40[48]=8'h60;
        mem_40[49]=8'h62;
        mem_40[50]=8'h64;
        mem_40[51]=8'h66;
        mem_40[52]=8'h68;
        mem_40[53]=8'h6a;
        mem_40[54]=8'h6c;
        mem_40[55]=8'h6e;
        mem_40[56]=8'h70;
        mem_40[57]=8'h72;
        mem_40[58]=8'h74;
        mem_40[59]=8'h76;
        mem_40[60]=8'h78;
        mem_40[61]=8'h7a;
        mem_40[62]=8'h7c;
        mem_40[63]=8'h7e;
        mem_40[64]=8'h80;
        mem_40[65]=8'h82;
        mem_40[66]=8'h84;
        mem_40[67]=8'h86;
        mem_40[68]=8'h88;
        mem_40[69]=8'h8a;
        mem_40[70]=8'h8c;
        mem_40[71]=8'h8e;
        mem_40[72]=8'h90;
        mem_40[73]=8'h92;
        mem_40[74]=8'h94;
        mem_40[75]=8'h96;
        mem_40[76]=8'h98;
        mem_40[77]=8'h9a;
        mem_40[78]=8'h9c;
        mem_40[79]=8'h9e;
        mem_40[80]=8'ha0;
        mem_40[81]=8'ha2;
        mem_40[82]=8'ha4;
        mem_40[83]=8'ha6;
        mem_40[84]=8'ha8;
        mem_40[85]=8'haa;
        mem_40[86]=8'hac;
        mem_40[87]=8'hae;
        mem_40[88]=8'hb0;
        mem_40[89]=8'hb2;
        mem_40[90]=8'hb4;
        mem_40[91]=8'hb6;
        mem_40[92]=8'hb8;
        mem_40[93]=8'hba;
        mem_40[94]=8'hbc;
        mem_40[95]=8'hbe;
        mem_40[96]=8'hc0;
        mem_40[97]=8'hc2;
        mem_40[98]=8'hc4;
        mem_40[99]=8'hc6;
        mem_40[100]=8'hc8;
        mem_40[101]=8'hca;
        mem_40[102]=8'hcc;
        mem_40[103]=8'hce;
        mem_40[104]=8'hd0;
        mem_40[105]=8'hd2;
        mem_40[106]=8'hd4;
        mem_40[107]=8'hd6;
        mem_40[108]=8'hd8;
        mem_40[109]=8'hda;
        mem_40[110]=8'hdc;
        mem_40[111]=8'hde;
        mem_40[112]=8'he0;
        mem_40[113]=8'he2;
        mem_40[114]=8'he4;
        mem_40[115]=8'he6;
        mem_40[116]=8'he8;
        mem_40[117]=8'hea;
        mem_40[118]=8'hec;
        mem_40[119]=8'hee;
        mem_40[120]=8'hf0;
        mem_40[121]=8'hf2;
        mem_40[122]=8'hf4;
        mem_40[123]=8'hf6;
        mem_40[124]=8'hf8;
        mem_40[125]=8'hfa;
        mem_40[126]=8'hfc;
        mem_40[127]=8'hfe;
        mem_40[128]=8'h1b;
        mem_40[129]=8'h19;
        mem_40[130]=8'h1f;
        mem_40[131]=8'h1d;
        mem_40[132]=8'h13;
        mem_40[133]=8'h11;
        mem_40[134]=8'h17;
        mem_40[135]=8'h15;
        mem_40[136]=8'hb;
        mem_40[137]=8'h9;
        mem_40[138]=8'hf;
        mem_40[139]=8'hd;
        mem_40[140]=8'h3;
        mem_40[141]=8'h1;
        mem_40[142]=8'h7;
        mem_40[143]=8'h5;
        mem_40[144]=8'h3b;
        mem_40[145]=8'h39;
        mem_40[146]=8'h3f;
        mem_40[147]=8'h3d;
        mem_40[148]=8'h33;
        mem_40[149]=8'h31;
        mem_40[150]=8'h37;
        mem_40[151]=8'h35;
        mem_40[152]=8'h2b;
        mem_40[153]=8'h29;
        mem_40[154]=8'h2f;
        mem_40[155]=8'h2d;
        mem_40[156]=8'h23;
        mem_40[157]=8'h21;
        mem_40[158]=8'h27;
        mem_40[159]=8'h25;
        mem_40[160]=8'h5b;
        mem_40[161]=8'h59;
        mem_40[162]=8'h5f;
        mem_40[163]=8'h5d;
        mem_40[164]=8'h53;
        mem_40[165]=8'h51;
        mem_40[166]=8'h57;
        mem_40[167]=8'h55;
        mem_40[168]=8'h4b;
        mem_40[169]=8'h49;
        mem_40[170]=8'h4f;
        mem_40[171]=8'h4d;
        mem_40[172]=8'h43;
        mem_40[173]=8'h41;
        mem_40[174]=8'h47;
        mem_40[175]=8'h45;
        mem_40[176]=8'h7b;
        mem_40[177]=8'h79;
        mem_40[178]=8'h7f;
        mem_40[179]=8'h7d;
        mem_40[180]=8'h73;
        mem_40[181]=8'h71;
        mem_40[182]=8'h77;
        mem_40[183]=8'h75;
        mem_40[184]=8'h6b;
        mem_40[185]=8'h69;
        mem_40[186]=8'h6f;
        mem_40[187]=8'h6d;
        mem_40[188]=8'h63;
        mem_40[189]=8'h61;
        mem_40[190]=8'h67;
        mem_40[191]=8'h65;
        mem_40[192]=8'h9b;
        mem_40[193]=8'h99;
        mem_40[194]=8'h9f;
        mem_40[195]=8'h9d;
        mem_40[196]=8'h93;
        mem_40[197]=8'h91;
        mem_40[198]=8'h97;
        mem_40[199]=8'h95;
        mem_40[200]=8'h8b;
        mem_40[201]=8'h89;
        mem_40[202]=8'h8f;
        mem_40[203]=8'h8d;
        mem_40[204]=8'h83;
        mem_40[205]=8'h81;
        mem_40[206]=8'h87;
        mem_40[207]=8'h85;
        mem_40[208]=8'hbb;
        mem_40[209]=8'hb9;
        mem_40[210]=8'hbf;
        mem_40[211]=8'hbd;
        mem_40[212]=8'hb3;
        mem_40[213]=8'hb1;
        mem_40[214]=8'hb7;
        mem_40[215]=8'hb5;
        mem_40[216]=8'hab;
        mem_40[217]=8'ha9;
        mem_40[218]=8'haf;
        mem_40[219]=8'had;
        mem_40[220]=8'ha3;
        mem_40[221]=8'ha1;
        mem_40[222]=8'ha7;
        mem_40[223]=8'ha5;
        mem_40[224]=8'hdb;
        mem_40[225]=8'hd9;
        mem_40[226]=8'hdf;
        mem_40[227]=8'hdd;
        mem_40[228]=8'hd3;
        mem_40[229]=8'hd1;
        mem_40[230]=8'hd7;
        mem_40[231]=8'hd5;
        mem_40[232]=8'hcb;
        mem_40[233]=8'hc9;
        mem_40[234]=8'hcf;
        mem_40[235]=8'hcd;
        mem_40[236]=8'hc3;
        mem_40[237]=8'hc1;
        mem_40[238]=8'hc7;
        mem_40[239]=8'hc5;
        mem_40[240]=8'hfb;
        mem_40[241]=8'hf9;
        mem_40[242]=8'hff;
        mem_40[243]=8'hfd;
        mem_40[244]=8'hf3;
        mem_40[245]=8'hf1;
        mem_40[246]=8'hf7;
        mem_40[247]=8'hf5;
        mem_40[248]=8'heb;
        mem_40[249]=8'he9;
        mem_40[250]=8'hef;
        mem_40[251]=8'hed;
        mem_40[252]=8'he3;
        mem_40[253]=8'he1;
        mem_40[254]=8'he7;
        mem_40[255]=8'he5;
    end

    initial begin
        mem_41[0]=8'h0;
        mem_41[1]=8'h3;
        mem_41[2]=8'h6;
        mem_41[3]=8'h5;
        mem_41[4]=8'hc;
        mem_41[5]=8'hf;
        mem_41[6]=8'ha;
        mem_41[7]=8'h9;
        mem_41[8]=8'h18;
        mem_41[9]=8'h1b;
        mem_41[10]=8'h1e;
        mem_41[11]=8'h1d;
        mem_41[12]=8'h14;
        mem_41[13]=8'h17;
        mem_41[14]=8'h12;
        mem_41[15]=8'h11;
        mem_41[16]=8'h30;
        mem_41[17]=8'h33;
        mem_41[18]=8'h36;
        mem_41[19]=8'h35;
        mem_41[20]=8'h3c;
        mem_41[21]=8'h3f;
        mem_41[22]=8'h3a;
        mem_41[23]=8'h39;
        mem_41[24]=8'h28;
        mem_41[25]=8'h2b;
        mem_41[26]=8'h2e;
        mem_41[27]=8'h2d;
        mem_41[28]=8'h24;
        mem_41[29]=8'h27;
        mem_41[30]=8'h22;
        mem_41[31]=8'h21;
        mem_41[32]=8'h60;
        mem_41[33]=8'h63;
        mem_41[34]=8'h66;
        mem_41[35]=8'h65;
        mem_41[36]=8'h6c;
        mem_41[37]=8'h6f;
        mem_41[38]=8'h6a;
        mem_41[39]=8'h69;
        mem_41[40]=8'h78;
        mem_41[41]=8'h7b;
        mem_41[42]=8'h7e;
        mem_41[43]=8'h7d;
        mem_41[44]=8'h74;
        mem_41[45]=8'h77;
        mem_41[46]=8'h72;
        mem_41[47]=8'h71;
        mem_41[48]=8'h50;
        mem_41[49]=8'h53;
        mem_41[50]=8'h56;
        mem_41[51]=8'h55;
        mem_41[52]=8'h5c;
        mem_41[53]=8'h5f;
        mem_41[54]=8'h5a;
        mem_41[55]=8'h59;
        mem_41[56]=8'h48;
        mem_41[57]=8'h4b;
        mem_41[58]=8'h4e;
        mem_41[59]=8'h4d;
        mem_41[60]=8'h44;
        mem_41[61]=8'h47;
        mem_41[62]=8'h42;
        mem_41[63]=8'h41;
        mem_41[64]=8'hc0;
        mem_41[65]=8'hc3;
        mem_41[66]=8'hc6;
        mem_41[67]=8'hc5;
        mem_41[68]=8'hcc;
        mem_41[69]=8'hcf;
        mem_41[70]=8'hca;
        mem_41[71]=8'hc9;
        mem_41[72]=8'hd8;
        mem_41[73]=8'hdb;
        mem_41[74]=8'hde;
        mem_41[75]=8'hdd;
        mem_41[76]=8'hd4;
        mem_41[77]=8'hd7;
        mem_41[78]=8'hd2;
        mem_41[79]=8'hd1;
        mem_41[80]=8'hf0;
        mem_41[81]=8'hf3;
        mem_41[82]=8'hf6;
        mem_41[83]=8'hf5;
        mem_41[84]=8'hfc;
        mem_41[85]=8'hff;
        mem_41[86]=8'hfa;
        mem_41[87]=8'hf9;
        mem_41[88]=8'he8;
        mem_41[89]=8'heb;
        mem_41[90]=8'hee;
        mem_41[91]=8'hed;
        mem_41[92]=8'he4;
        mem_41[93]=8'he7;
        mem_41[94]=8'he2;
        mem_41[95]=8'he1;
        mem_41[96]=8'ha0;
        mem_41[97]=8'ha3;
        mem_41[98]=8'ha6;
        mem_41[99]=8'ha5;
        mem_41[100]=8'hac;
        mem_41[101]=8'haf;
        mem_41[102]=8'haa;
        mem_41[103]=8'ha9;
        mem_41[104]=8'hb8;
        mem_41[105]=8'hbb;
        mem_41[106]=8'hbe;
        mem_41[107]=8'hbd;
        mem_41[108]=8'hb4;
        mem_41[109]=8'hb7;
        mem_41[110]=8'hb2;
        mem_41[111]=8'hb1;
        mem_41[112]=8'h90;
        mem_41[113]=8'h93;
        mem_41[114]=8'h96;
        mem_41[115]=8'h95;
        mem_41[116]=8'h9c;
        mem_41[117]=8'h9f;
        mem_41[118]=8'h9a;
        mem_41[119]=8'h99;
        mem_41[120]=8'h88;
        mem_41[121]=8'h8b;
        mem_41[122]=8'h8e;
        mem_41[123]=8'h8d;
        mem_41[124]=8'h84;
        mem_41[125]=8'h87;
        mem_41[126]=8'h82;
        mem_41[127]=8'h81;
        mem_41[128]=8'h9b;
        mem_41[129]=8'h98;
        mem_41[130]=8'h9d;
        mem_41[131]=8'h9e;
        mem_41[132]=8'h97;
        mem_41[133]=8'h94;
        mem_41[134]=8'h91;
        mem_41[135]=8'h92;
        mem_41[136]=8'h83;
        mem_41[137]=8'h80;
        mem_41[138]=8'h85;
        mem_41[139]=8'h86;
        mem_41[140]=8'h8f;
        mem_41[141]=8'h8c;
        mem_41[142]=8'h89;
        mem_41[143]=8'h8a;
        mem_41[144]=8'hab;
        mem_41[145]=8'ha8;
        mem_41[146]=8'had;
        mem_41[147]=8'hae;
        mem_41[148]=8'ha7;
        mem_41[149]=8'ha4;
        mem_41[150]=8'ha1;
        mem_41[151]=8'ha2;
        mem_41[152]=8'hb3;
        mem_41[153]=8'hb0;
        mem_41[154]=8'hb5;
        mem_41[155]=8'hb6;
        mem_41[156]=8'hbf;
        mem_41[157]=8'hbc;
        mem_41[158]=8'hb9;
        mem_41[159]=8'hba;
        mem_41[160]=8'hfb;
        mem_41[161]=8'hf8;
        mem_41[162]=8'hfd;
        mem_41[163]=8'hfe;
        mem_41[164]=8'hf7;
        mem_41[165]=8'hf4;
        mem_41[166]=8'hf1;
        mem_41[167]=8'hf2;
        mem_41[168]=8'he3;
        mem_41[169]=8'he0;
        mem_41[170]=8'he5;
        mem_41[171]=8'he6;
        mem_41[172]=8'hef;
        mem_41[173]=8'hec;
        mem_41[174]=8'he9;
        mem_41[175]=8'hea;
        mem_41[176]=8'hcb;
        mem_41[177]=8'hc8;
        mem_41[178]=8'hcd;
        mem_41[179]=8'hce;
        mem_41[180]=8'hc7;
        mem_41[181]=8'hc4;
        mem_41[182]=8'hc1;
        mem_41[183]=8'hc2;
        mem_41[184]=8'hd3;
        mem_41[185]=8'hd0;
        mem_41[186]=8'hd5;
        mem_41[187]=8'hd6;
        mem_41[188]=8'hdf;
        mem_41[189]=8'hdc;
        mem_41[190]=8'hd9;
        mem_41[191]=8'hda;
        mem_41[192]=8'h5b;
        mem_41[193]=8'h58;
        mem_41[194]=8'h5d;
        mem_41[195]=8'h5e;
        mem_41[196]=8'h57;
        mem_41[197]=8'h54;
        mem_41[198]=8'h51;
        mem_41[199]=8'h52;
        mem_41[200]=8'h43;
        mem_41[201]=8'h40;
        mem_41[202]=8'h45;
        mem_41[203]=8'h46;
        mem_41[204]=8'h4f;
        mem_41[205]=8'h4c;
        mem_41[206]=8'h49;
        mem_41[207]=8'h4a;
        mem_41[208]=8'h6b;
        mem_41[209]=8'h68;
        mem_41[210]=8'h6d;
        mem_41[211]=8'h6e;
        mem_41[212]=8'h67;
        mem_41[213]=8'h64;
        mem_41[214]=8'h61;
        mem_41[215]=8'h62;
        mem_41[216]=8'h73;
        mem_41[217]=8'h70;
        mem_41[218]=8'h75;
        mem_41[219]=8'h76;
        mem_41[220]=8'h7f;
        mem_41[221]=8'h7c;
        mem_41[222]=8'h79;
        mem_41[223]=8'h7a;
        mem_41[224]=8'h3b;
        mem_41[225]=8'h38;
        mem_41[226]=8'h3d;
        mem_41[227]=8'h3e;
        mem_41[228]=8'h37;
        mem_41[229]=8'h34;
        mem_41[230]=8'h31;
        mem_41[231]=8'h32;
        mem_41[232]=8'h23;
        mem_41[233]=8'h20;
        mem_41[234]=8'h25;
        mem_41[235]=8'h26;
        mem_41[236]=8'h2f;
        mem_41[237]=8'h2c;
        mem_41[238]=8'h29;
        mem_41[239]=8'h2a;
        mem_41[240]=8'hb;
        mem_41[241]=8'h8;
        mem_41[242]=8'hd;
        mem_41[243]=8'he;
        mem_41[244]=8'h7;
        mem_41[245]=8'h4;
        mem_41[246]=8'h1;
        mem_41[247]=8'h2;
        mem_41[248]=8'h13;
        mem_41[249]=8'h10;
        mem_41[250]=8'h15;
        mem_41[251]=8'h16;
        mem_41[252]=8'h1f;
        mem_41[253]=8'h1c;
        mem_41[254]=8'h19;
        mem_41[255]=8'h1a;
    end

    initial begin
        mem_42[0]=8'h0;
        mem_42[1]=8'h2;
        mem_42[2]=8'h4;
        mem_42[3]=8'h6;
        mem_42[4]=8'h8;
        mem_42[5]=8'ha;
        mem_42[6]=8'hc;
        mem_42[7]=8'he;
        mem_42[8]=8'h10;
        mem_42[9]=8'h12;
        mem_42[10]=8'h14;
        mem_42[11]=8'h16;
        mem_42[12]=8'h18;
        mem_42[13]=8'h1a;
        mem_42[14]=8'h1c;
        mem_42[15]=8'h1e;
        mem_42[16]=8'h20;
        mem_42[17]=8'h22;
        mem_42[18]=8'h24;
        mem_42[19]=8'h26;
        mem_42[20]=8'h28;
        mem_42[21]=8'h2a;
        mem_42[22]=8'h2c;
        mem_42[23]=8'h2e;
        mem_42[24]=8'h30;
        mem_42[25]=8'h32;
        mem_42[26]=8'h34;
        mem_42[27]=8'h36;
        mem_42[28]=8'h38;
        mem_42[29]=8'h3a;
        mem_42[30]=8'h3c;
        mem_42[31]=8'h3e;
        mem_42[32]=8'h40;
        mem_42[33]=8'h42;
        mem_42[34]=8'h44;
        mem_42[35]=8'h46;
        mem_42[36]=8'h48;
        mem_42[37]=8'h4a;
        mem_42[38]=8'h4c;
        mem_42[39]=8'h4e;
        mem_42[40]=8'h50;
        mem_42[41]=8'h52;
        mem_42[42]=8'h54;
        mem_42[43]=8'h56;
        mem_42[44]=8'h58;
        mem_42[45]=8'h5a;
        mem_42[46]=8'h5c;
        mem_42[47]=8'h5e;
        mem_42[48]=8'h60;
        mem_42[49]=8'h62;
        mem_42[50]=8'h64;
        mem_42[51]=8'h66;
        mem_42[52]=8'h68;
        mem_42[53]=8'h6a;
        mem_42[54]=8'h6c;
        mem_42[55]=8'h6e;
        mem_42[56]=8'h70;
        mem_42[57]=8'h72;
        mem_42[58]=8'h74;
        mem_42[59]=8'h76;
        mem_42[60]=8'h78;
        mem_42[61]=8'h7a;
        mem_42[62]=8'h7c;
        mem_42[63]=8'h7e;
        mem_42[64]=8'h80;
        mem_42[65]=8'h82;
        mem_42[66]=8'h84;
        mem_42[67]=8'h86;
        mem_42[68]=8'h88;
        mem_42[69]=8'h8a;
        mem_42[70]=8'h8c;
        mem_42[71]=8'h8e;
        mem_42[72]=8'h90;
        mem_42[73]=8'h92;
        mem_42[74]=8'h94;
        mem_42[75]=8'h96;
        mem_42[76]=8'h98;
        mem_42[77]=8'h9a;
        mem_42[78]=8'h9c;
        mem_42[79]=8'h9e;
        mem_42[80]=8'ha0;
        mem_42[81]=8'ha2;
        mem_42[82]=8'ha4;
        mem_42[83]=8'ha6;
        mem_42[84]=8'ha8;
        mem_42[85]=8'haa;
        mem_42[86]=8'hac;
        mem_42[87]=8'hae;
        mem_42[88]=8'hb0;
        mem_42[89]=8'hb2;
        mem_42[90]=8'hb4;
        mem_42[91]=8'hb6;
        mem_42[92]=8'hb8;
        mem_42[93]=8'hba;
        mem_42[94]=8'hbc;
        mem_42[95]=8'hbe;
        mem_42[96]=8'hc0;
        mem_42[97]=8'hc2;
        mem_42[98]=8'hc4;
        mem_42[99]=8'hc6;
        mem_42[100]=8'hc8;
        mem_42[101]=8'hca;
        mem_42[102]=8'hcc;
        mem_42[103]=8'hce;
        mem_42[104]=8'hd0;
        mem_42[105]=8'hd2;
        mem_42[106]=8'hd4;
        mem_42[107]=8'hd6;
        mem_42[108]=8'hd8;
        mem_42[109]=8'hda;
        mem_42[110]=8'hdc;
        mem_42[111]=8'hde;
        mem_42[112]=8'he0;
        mem_42[113]=8'he2;
        mem_42[114]=8'he4;
        mem_42[115]=8'he6;
        mem_42[116]=8'he8;
        mem_42[117]=8'hea;
        mem_42[118]=8'hec;
        mem_42[119]=8'hee;
        mem_42[120]=8'hf0;
        mem_42[121]=8'hf2;
        mem_42[122]=8'hf4;
        mem_42[123]=8'hf6;
        mem_42[124]=8'hf8;
        mem_42[125]=8'hfa;
        mem_42[126]=8'hfc;
        mem_42[127]=8'hfe;
        mem_42[128]=8'h1b;
        mem_42[129]=8'h19;
        mem_42[130]=8'h1f;
        mem_42[131]=8'h1d;
        mem_42[132]=8'h13;
        mem_42[133]=8'h11;
        mem_42[134]=8'h17;
        mem_42[135]=8'h15;
        mem_42[136]=8'hb;
        mem_42[137]=8'h9;
        mem_42[138]=8'hf;
        mem_42[139]=8'hd;
        mem_42[140]=8'h3;
        mem_42[141]=8'h1;
        mem_42[142]=8'h7;
        mem_42[143]=8'h5;
        mem_42[144]=8'h3b;
        mem_42[145]=8'h39;
        mem_42[146]=8'h3f;
        mem_42[147]=8'h3d;
        mem_42[148]=8'h33;
        mem_42[149]=8'h31;
        mem_42[150]=8'h37;
        mem_42[151]=8'h35;
        mem_42[152]=8'h2b;
        mem_42[153]=8'h29;
        mem_42[154]=8'h2f;
        mem_42[155]=8'h2d;
        mem_42[156]=8'h23;
        mem_42[157]=8'h21;
        mem_42[158]=8'h27;
        mem_42[159]=8'h25;
        mem_42[160]=8'h5b;
        mem_42[161]=8'h59;
        mem_42[162]=8'h5f;
        mem_42[163]=8'h5d;
        mem_42[164]=8'h53;
        mem_42[165]=8'h51;
        mem_42[166]=8'h57;
        mem_42[167]=8'h55;
        mem_42[168]=8'h4b;
        mem_42[169]=8'h49;
        mem_42[170]=8'h4f;
        mem_42[171]=8'h4d;
        mem_42[172]=8'h43;
        mem_42[173]=8'h41;
        mem_42[174]=8'h47;
        mem_42[175]=8'h45;
        mem_42[176]=8'h7b;
        mem_42[177]=8'h79;
        mem_42[178]=8'h7f;
        mem_42[179]=8'h7d;
        mem_42[180]=8'h73;
        mem_42[181]=8'h71;
        mem_42[182]=8'h77;
        mem_42[183]=8'h75;
        mem_42[184]=8'h6b;
        mem_42[185]=8'h69;
        mem_42[186]=8'h6f;
        mem_42[187]=8'h6d;
        mem_42[188]=8'h63;
        mem_42[189]=8'h61;
        mem_42[190]=8'h67;
        mem_42[191]=8'h65;
        mem_42[192]=8'h9b;
        mem_42[193]=8'h99;
        mem_42[194]=8'h9f;
        mem_42[195]=8'h9d;
        mem_42[196]=8'h93;
        mem_42[197]=8'h91;
        mem_42[198]=8'h97;
        mem_42[199]=8'h95;
        mem_42[200]=8'h8b;
        mem_42[201]=8'h89;
        mem_42[202]=8'h8f;
        mem_42[203]=8'h8d;
        mem_42[204]=8'h83;
        mem_42[205]=8'h81;
        mem_42[206]=8'h87;
        mem_42[207]=8'h85;
        mem_42[208]=8'hbb;
        mem_42[209]=8'hb9;
        mem_42[210]=8'hbf;
        mem_42[211]=8'hbd;
        mem_42[212]=8'hb3;
        mem_42[213]=8'hb1;
        mem_42[214]=8'hb7;
        mem_42[215]=8'hb5;
        mem_42[216]=8'hab;
        mem_42[217]=8'ha9;
        mem_42[218]=8'haf;
        mem_42[219]=8'had;
        mem_42[220]=8'ha3;
        mem_42[221]=8'ha1;
        mem_42[222]=8'ha7;
        mem_42[223]=8'ha5;
        mem_42[224]=8'hdb;
        mem_42[225]=8'hd9;
        mem_42[226]=8'hdf;
        mem_42[227]=8'hdd;
        mem_42[228]=8'hd3;
        mem_42[229]=8'hd1;
        mem_42[230]=8'hd7;
        mem_42[231]=8'hd5;
        mem_42[232]=8'hcb;
        mem_42[233]=8'hc9;
        mem_42[234]=8'hcf;
        mem_42[235]=8'hcd;
        mem_42[236]=8'hc3;
        mem_42[237]=8'hc1;
        mem_42[238]=8'hc7;
        mem_42[239]=8'hc5;
        mem_42[240]=8'hfb;
        mem_42[241]=8'hf9;
        mem_42[242]=8'hff;
        mem_42[243]=8'hfd;
        mem_42[244]=8'hf3;
        mem_42[245]=8'hf1;
        mem_42[246]=8'hf7;
        mem_42[247]=8'hf5;
        mem_42[248]=8'heb;
        mem_42[249]=8'he9;
        mem_42[250]=8'hef;
        mem_42[251]=8'hed;
        mem_42[252]=8'he3;
        mem_42[253]=8'he1;
        mem_42[254]=8'he7;
        mem_42[255]=8'he5;
    end

    initial begin
        mem_43[0]=8'h0;
        mem_43[1]=8'h3;
        mem_43[2]=8'h6;
        mem_43[3]=8'h5;
        mem_43[4]=8'hc;
        mem_43[5]=8'hf;
        mem_43[6]=8'ha;
        mem_43[7]=8'h9;
        mem_43[8]=8'h18;
        mem_43[9]=8'h1b;
        mem_43[10]=8'h1e;
        mem_43[11]=8'h1d;
        mem_43[12]=8'h14;
        mem_43[13]=8'h17;
        mem_43[14]=8'h12;
        mem_43[15]=8'h11;
        mem_43[16]=8'h30;
        mem_43[17]=8'h33;
        mem_43[18]=8'h36;
        mem_43[19]=8'h35;
        mem_43[20]=8'h3c;
        mem_43[21]=8'h3f;
        mem_43[22]=8'h3a;
        mem_43[23]=8'h39;
        mem_43[24]=8'h28;
        mem_43[25]=8'h2b;
        mem_43[26]=8'h2e;
        mem_43[27]=8'h2d;
        mem_43[28]=8'h24;
        mem_43[29]=8'h27;
        mem_43[30]=8'h22;
        mem_43[31]=8'h21;
        mem_43[32]=8'h60;
        mem_43[33]=8'h63;
        mem_43[34]=8'h66;
        mem_43[35]=8'h65;
        mem_43[36]=8'h6c;
        mem_43[37]=8'h6f;
        mem_43[38]=8'h6a;
        mem_43[39]=8'h69;
        mem_43[40]=8'h78;
        mem_43[41]=8'h7b;
        mem_43[42]=8'h7e;
        mem_43[43]=8'h7d;
        mem_43[44]=8'h74;
        mem_43[45]=8'h77;
        mem_43[46]=8'h72;
        mem_43[47]=8'h71;
        mem_43[48]=8'h50;
        mem_43[49]=8'h53;
        mem_43[50]=8'h56;
        mem_43[51]=8'h55;
        mem_43[52]=8'h5c;
        mem_43[53]=8'h5f;
        mem_43[54]=8'h5a;
        mem_43[55]=8'h59;
        mem_43[56]=8'h48;
        mem_43[57]=8'h4b;
        mem_43[58]=8'h4e;
        mem_43[59]=8'h4d;
        mem_43[60]=8'h44;
        mem_43[61]=8'h47;
        mem_43[62]=8'h42;
        mem_43[63]=8'h41;
        mem_43[64]=8'hc0;
        mem_43[65]=8'hc3;
        mem_43[66]=8'hc6;
        mem_43[67]=8'hc5;
        mem_43[68]=8'hcc;
        mem_43[69]=8'hcf;
        mem_43[70]=8'hca;
        mem_43[71]=8'hc9;
        mem_43[72]=8'hd8;
        mem_43[73]=8'hdb;
        mem_43[74]=8'hde;
        mem_43[75]=8'hdd;
        mem_43[76]=8'hd4;
        mem_43[77]=8'hd7;
        mem_43[78]=8'hd2;
        mem_43[79]=8'hd1;
        mem_43[80]=8'hf0;
        mem_43[81]=8'hf3;
        mem_43[82]=8'hf6;
        mem_43[83]=8'hf5;
        mem_43[84]=8'hfc;
        mem_43[85]=8'hff;
        mem_43[86]=8'hfa;
        mem_43[87]=8'hf9;
        mem_43[88]=8'he8;
        mem_43[89]=8'heb;
        mem_43[90]=8'hee;
        mem_43[91]=8'hed;
        mem_43[92]=8'he4;
        mem_43[93]=8'he7;
        mem_43[94]=8'he2;
        mem_43[95]=8'he1;
        mem_43[96]=8'ha0;
        mem_43[97]=8'ha3;
        mem_43[98]=8'ha6;
        mem_43[99]=8'ha5;
        mem_43[100]=8'hac;
        mem_43[101]=8'haf;
        mem_43[102]=8'haa;
        mem_43[103]=8'ha9;
        mem_43[104]=8'hb8;
        mem_43[105]=8'hbb;
        mem_43[106]=8'hbe;
        mem_43[107]=8'hbd;
        mem_43[108]=8'hb4;
        mem_43[109]=8'hb7;
        mem_43[110]=8'hb2;
        mem_43[111]=8'hb1;
        mem_43[112]=8'h90;
        mem_43[113]=8'h93;
        mem_43[114]=8'h96;
        mem_43[115]=8'h95;
        mem_43[116]=8'h9c;
        mem_43[117]=8'h9f;
        mem_43[118]=8'h9a;
        mem_43[119]=8'h99;
        mem_43[120]=8'h88;
        mem_43[121]=8'h8b;
        mem_43[122]=8'h8e;
        mem_43[123]=8'h8d;
        mem_43[124]=8'h84;
        mem_43[125]=8'h87;
        mem_43[126]=8'h82;
        mem_43[127]=8'h81;
        mem_43[128]=8'h9b;
        mem_43[129]=8'h98;
        mem_43[130]=8'h9d;
        mem_43[131]=8'h9e;
        mem_43[132]=8'h97;
        mem_43[133]=8'h94;
        mem_43[134]=8'h91;
        mem_43[135]=8'h92;
        mem_43[136]=8'h83;
        mem_43[137]=8'h80;
        mem_43[138]=8'h85;
        mem_43[139]=8'h86;
        mem_43[140]=8'h8f;
        mem_43[141]=8'h8c;
        mem_43[142]=8'h89;
        mem_43[143]=8'h8a;
        mem_43[144]=8'hab;
        mem_43[145]=8'ha8;
        mem_43[146]=8'had;
        mem_43[147]=8'hae;
        mem_43[148]=8'ha7;
        mem_43[149]=8'ha4;
        mem_43[150]=8'ha1;
        mem_43[151]=8'ha2;
        mem_43[152]=8'hb3;
        mem_43[153]=8'hb0;
        mem_43[154]=8'hb5;
        mem_43[155]=8'hb6;
        mem_43[156]=8'hbf;
        mem_43[157]=8'hbc;
        mem_43[158]=8'hb9;
        mem_43[159]=8'hba;
        mem_43[160]=8'hfb;
        mem_43[161]=8'hf8;
        mem_43[162]=8'hfd;
        mem_43[163]=8'hfe;
        mem_43[164]=8'hf7;
        mem_43[165]=8'hf4;
        mem_43[166]=8'hf1;
        mem_43[167]=8'hf2;
        mem_43[168]=8'he3;
        mem_43[169]=8'he0;
        mem_43[170]=8'he5;
        mem_43[171]=8'he6;
        mem_43[172]=8'hef;
        mem_43[173]=8'hec;
        mem_43[174]=8'he9;
        mem_43[175]=8'hea;
        mem_43[176]=8'hcb;
        mem_43[177]=8'hc8;
        mem_43[178]=8'hcd;
        mem_43[179]=8'hce;
        mem_43[180]=8'hc7;
        mem_43[181]=8'hc4;
        mem_43[182]=8'hc1;
        mem_43[183]=8'hc2;
        mem_43[184]=8'hd3;
        mem_43[185]=8'hd0;
        mem_43[186]=8'hd5;
        mem_43[187]=8'hd6;
        mem_43[188]=8'hdf;
        mem_43[189]=8'hdc;
        mem_43[190]=8'hd9;
        mem_43[191]=8'hda;
        mem_43[192]=8'h5b;
        mem_43[193]=8'h58;
        mem_43[194]=8'h5d;
        mem_43[195]=8'h5e;
        mem_43[196]=8'h57;
        mem_43[197]=8'h54;
        mem_43[198]=8'h51;
        mem_43[199]=8'h52;
        mem_43[200]=8'h43;
        mem_43[201]=8'h40;
        mem_43[202]=8'h45;
        mem_43[203]=8'h46;
        mem_43[204]=8'h4f;
        mem_43[205]=8'h4c;
        mem_43[206]=8'h49;
        mem_43[207]=8'h4a;
        mem_43[208]=8'h6b;
        mem_43[209]=8'h68;
        mem_43[210]=8'h6d;
        mem_43[211]=8'h6e;
        mem_43[212]=8'h67;
        mem_43[213]=8'h64;
        mem_43[214]=8'h61;
        mem_43[215]=8'h62;
        mem_43[216]=8'h73;
        mem_43[217]=8'h70;
        mem_43[218]=8'h75;
        mem_43[219]=8'h76;
        mem_43[220]=8'h7f;
        mem_43[221]=8'h7c;
        mem_43[222]=8'h79;
        mem_43[223]=8'h7a;
        mem_43[224]=8'h3b;
        mem_43[225]=8'h38;
        mem_43[226]=8'h3d;
        mem_43[227]=8'h3e;
        mem_43[228]=8'h37;
        mem_43[229]=8'h34;
        mem_43[230]=8'h31;
        mem_43[231]=8'h32;
        mem_43[232]=8'h23;
        mem_43[233]=8'h20;
        mem_43[234]=8'h25;
        mem_43[235]=8'h26;
        mem_43[236]=8'h2f;
        mem_43[237]=8'h2c;
        mem_43[238]=8'h29;
        mem_43[239]=8'h2a;
        mem_43[240]=8'hb;
        mem_43[241]=8'h8;
        mem_43[242]=8'hd;
        mem_43[243]=8'he;
        mem_43[244]=8'h7;
        mem_43[245]=8'h4;
        mem_43[246]=8'h1;
        mem_43[247]=8'h2;
        mem_43[248]=8'h13;
        mem_43[249]=8'h10;
        mem_43[250]=8'h15;
        mem_43[251]=8'h16;
        mem_43[252]=8'h1f;
        mem_43[253]=8'h1c;
        mem_43[254]=8'h19;
        mem_43[255]=8'h1a;
    end

    initial begin
        mem_44[0]=8'h0;
        mem_44[1]=8'h2;
        mem_44[2]=8'h4;
        mem_44[3]=8'h6;
        mem_44[4]=8'h8;
        mem_44[5]=8'ha;
        mem_44[6]=8'hc;
        mem_44[7]=8'he;
        mem_44[8]=8'h10;
        mem_44[9]=8'h12;
        mem_44[10]=8'h14;
        mem_44[11]=8'h16;
        mem_44[12]=8'h18;
        mem_44[13]=8'h1a;
        mem_44[14]=8'h1c;
        mem_44[15]=8'h1e;
        mem_44[16]=8'h20;
        mem_44[17]=8'h22;
        mem_44[18]=8'h24;
        mem_44[19]=8'h26;
        mem_44[20]=8'h28;
        mem_44[21]=8'h2a;
        mem_44[22]=8'h2c;
        mem_44[23]=8'h2e;
        mem_44[24]=8'h30;
        mem_44[25]=8'h32;
        mem_44[26]=8'h34;
        mem_44[27]=8'h36;
        mem_44[28]=8'h38;
        mem_44[29]=8'h3a;
        mem_44[30]=8'h3c;
        mem_44[31]=8'h3e;
        mem_44[32]=8'h40;
        mem_44[33]=8'h42;
        mem_44[34]=8'h44;
        mem_44[35]=8'h46;
        mem_44[36]=8'h48;
        mem_44[37]=8'h4a;
        mem_44[38]=8'h4c;
        mem_44[39]=8'h4e;
        mem_44[40]=8'h50;
        mem_44[41]=8'h52;
        mem_44[42]=8'h54;
        mem_44[43]=8'h56;
        mem_44[44]=8'h58;
        mem_44[45]=8'h5a;
        mem_44[46]=8'h5c;
        mem_44[47]=8'h5e;
        mem_44[48]=8'h60;
        mem_44[49]=8'h62;
        mem_44[50]=8'h64;
        mem_44[51]=8'h66;
        mem_44[52]=8'h68;
        mem_44[53]=8'h6a;
        mem_44[54]=8'h6c;
        mem_44[55]=8'h6e;
        mem_44[56]=8'h70;
        mem_44[57]=8'h72;
        mem_44[58]=8'h74;
        mem_44[59]=8'h76;
        mem_44[60]=8'h78;
        mem_44[61]=8'h7a;
        mem_44[62]=8'h7c;
        mem_44[63]=8'h7e;
        mem_44[64]=8'h80;
        mem_44[65]=8'h82;
        mem_44[66]=8'h84;
        mem_44[67]=8'h86;
        mem_44[68]=8'h88;
        mem_44[69]=8'h8a;
        mem_44[70]=8'h8c;
        mem_44[71]=8'h8e;
        mem_44[72]=8'h90;
        mem_44[73]=8'h92;
        mem_44[74]=8'h94;
        mem_44[75]=8'h96;
        mem_44[76]=8'h98;
        mem_44[77]=8'h9a;
        mem_44[78]=8'h9c;
        mem_44[79]=8'h9e;
        mem_44[80]=8'ha0;
        mem_44[81]=8'ha2;
        mem_44[82]=8'ha4;
        mem_44[83]=8'ha6;
        mem_44[84]=8'ha8;
        mem_44[85]=8'haa;
        mem_44[86]=8'hac;
        mem_44[87]=8'hae;
        mem_44[88]=8'hb0;
        mem_44[89]=8'hb2;
        mem_44[90]=8'hb4;
        mem_44[91]=8'hb6;
        mem_44[92]=8'hb8;
        mem_44[93]=8'hba;
        mem_44[94]=8'hbc;
        mem_44[95]=8'hbe;
        mem_44[96]=8'hc0;
        mem_44[97]=8'hc2;
        mem_44[98]=8'hc4;
        mem_44[99]=8'hc6;
        mem_44[100]=8'hc8;
        mem_44[101]=8'hca;
        mem_44[102]=8'hcc;
        mem_44[103]=8'hce;
        mem_44[104]=8'hd0;
        mem_44[105]=8'hd2;
        mem_44[106]=8'hd4;
        mem_44[107]=8'hd6;
        mem_44[108]=8'hd8;
        mem_44[109]=8'hda;
        mem_44[110]=8'hdc;
        mem_44[111]=8'hde;
        mem_44[112]=8'he0;
        mem_44[113]=8'he2;
        mem_44[114]=8'he4;
        mem_44[115]=8'he6;
        mem_44[116]=8'he8;
        mem_44[117]=8'hea;
        mem_44[118]=8'hec;
        mem_44[119]=8'hee;
        mem_44[120]=8'hf0;
        mem_44[121]=8'hf2;
        mem_44[122]=8'hf4;
        mem_44[123]=8'hf6;
        mem_44[124]=8'hf8;
        mem_44[125]=8'hfa;
        mem_44[126]=8'hfc;
        mem_44[127]=8'hfe;
        mem_44[128]=8'h1b;
        mem_44[129]=8'h19;
        mem_44[130]=8'h1f;
        mem_44[131]=8'h1d;
        mem_44[132]=8'h13;
        mem_44[133]=8'h11;
        mem_44[134]=8'h17;
        mem_44[135]=8'h15;
        mem_44[136]=8'hb;
        mem_44[137]=8'h9;
        mem_44[138]=8'hf;
        mem_44[139]=8'hd;
        mem_44[140]=8'h3;
        mem_44[141]=8'h1;
        mem_44[142]=8'h7;
        mem_44[143]=8'h5;
        mem_44[144]=8'h3b;
        mem_44[145]=8'h39;
        mem_44[146]=8'h3f;
        mem_44[147]=8'h3d;
        mem_44[148]=8'h33;
        mem_44[149]=8'h31;
        mem_44[150]=8'h37;
        mem_44[151]=8'h35;
        mem_44[152]=8'h2b;
        mem_44[153]=8'h29;
        mem_44[154]=8'h2f;
        mem_44[155]=8'h2d;
        mem_44[156]=8'h23;
        mem_44[157]=8'h21;
        mem_44[158]=8'h27;
        mem_44[159]=8'h25;
        mem_44[160]=8'h5b;
        mem_44[161]=8'h59;
        mem_44[162]=8'h5f;
        mem_44[163]=8'h5d;
        mem_44[164]=8'h53;
        mem_44[165]=8'h51;
        mem_44[166]=8'h57;
        mem_44[167]=8'h55;
        mem_44[168]=8'h4b;
        mem_44[169]=8'h49;
        mem_44[170]=8'h4f;
        mem_44[171]=8'h4d;
        mem_44[172]=8'h43;
        mem_44[173]=8'h41;
        mem_44[174]=8'h47;
        mem_44[175]=8'h45;
        mem_44[176]=8'h7b;
        mem_44[177]=8'h79;
        mem_44[178]=8'h7f;
        mem_44[179]=8'h7d;
        mem_44[180]=8'h73;
        mem_44[181]=8'h71;
        mem_44[182]=8'h77;
        mem_44[183]=8'h75;
        mem_44[184]=8'h6b;
        mem_44[185]=8'h69;
        mem_44[186]=8'h6f;
        mem_44[187]=8'h6d;
        mem_44[188]=8'h63;
        mem_44[189]=8'h61;
        mem_44[190]=8'h67;
        mem_44[191]=8'h65;
        mem_44[192]=8'h9b;
        mem_44[193]=8'h99;
        mem_44[194]=8'h9f;
        mem_44[195]=8'h9d;
        mem_44[196]=8'h93;
        mem_44[197]=8'h91;
        mem_44[198]=8'h97;
        mem_44[199]=8'h95;
        mem_44[200]=8'h8b;
        mem_44[201]=8'h89;
        mem_44[202]=8'h8f;
        mem_44[203]=8'h8d;
        mem_44[204]=8'h83;
        mem_44[205]=8'h81;
        mem_44[206]=8'h87;
        mem_44[207]=8'h85;
        mem_44[208]=8'hbb;
        mem_44[209]=8'hb9;
        mem_44[210]=8'hbf;
        mem_44[211]=8'hbd;
        mem_44[212]=8'hb3;
        mem_44[213]=8'hb1;
        mem_44[214]=8'hb7;
        mem_44[215]=8'hb5;
        mem_44[216]=8'hab;
        mem_44[217]=8'ha9;
        mem_44[218]=8'haf;
        mem_44[219]=8'had;
        mem_44[220]=8'ha3;
        mem_44[221]=8'ha1;
        mem_44[222]=8'ha7;
        mem_44[223]=8'ha5;
        mem_44[224]=8'hdb;
        mem_44[225]=8'hd9;
        mem_44[226]=8'hdf;
        mem_44[227]=8'hdd;
        mem_44[228]=8'hd3;
        mem_44[229]=8'hd1;
        mem_44[230]=8'hd7;
        mem_44[231]=8'hd5;
        mem_44[232]=8'hcb;
        mem_44[233]=8'hc9;
        mem_44[234]=8'hcf;
        mem_44[235]=8'hcd;
        mem_44[236]=8'hc3;
        mem_44[237]=8'hc1;
        mem_44[238]=8'hc7;
        mem_44[239]=8'hc5;
        mem_44[240]=8'hfb;
        mem_44[241]=8'hf9;
        mem_44[242]=8'hff;
        mem_44[243]=8'hfd;
        mem_44[244]=8'hf3;
        mem_44[245]=8'hf1;
        mem_44[246]=8'hf7;
        mem_44[247]=8'hf5;
        mem_44[248]=8'heb;
        mem_44[249]=8'he9;
        mem_44[250]=8'hef;
        mem_44[251]=8'hed;
        mem_44[252]=8'he3;
        mem_44[253]=8'he1;
        mem_44[254]=8'he7;
        mem_44[255]=8'he5;
    end

    initial begin
        mem_45[0]=8'h0;
        mem_45[1]=8'h3;
        mem_45[2]=8'h6;
        mem_45[3]=8'h5;
        mem_45[4]=8'hc;
        mem_45[5]=8'hf;
        mem_45[6]=8'ha;
        mem_45[7]=8'h9;
        mem_45[8]=8'h18;
        mem_45[9]=8'h1b;
        mem_45[10]=8'h1e;
        mem_45[11]=8'h1d;
        mem_45[12]=8'h14;
        mem_45[13]=8'h17;
        mem_45[14]=8'h12;
        mem_45[15]=8'h11;
        mem_45[16]=8'h30;
        mem_45[17]=8'h33;
        mem_45[18]=8'h36;
        mem_45[19]=8'h35;
        mem_45[20]=8'h3c;
        mem_45[21]=8'h3f;
        mem_45[22]=8'h3a;
        mem_45[23]=8'h39;
        mem_45[24]=8'h28;
        mem_45[25]=8'h2b;
        mem_45[26]=8'h2e;
        mem_45[27]=8'h2d;
        mem_45[28]=8'h24;
        mem_45[29]=8'h27;
        mem_45[30]=8'h22;
        mem_45[31]=8'h21;
        mem_45[32]=8'h60;
        mem_45[33]=8'h63;
        mem_45[34]=8'h66;
        mem_45[35]=8'h65;
        mem_45[36]=8'h6c;
        mem_45[37]=8'h6f;
        mem_45[38]=8'h6a;
        mem_45[39]=8'h69;
        mem_45[40]=8'h78;
        mem_45[41]=8'h7b;
        mem_45[42]=8'h7e;
        mem_45[43]=8'h7d;
        mem_45[44]=8'h74;
        mem_45[45]=8'h77;
        mem_45[46]=8'h72;
        mem_45[47]=8'h71;
        mem_45[48]=8'h50;
        mem_45[49]=8'h53;
        mem_45[50]=8'h56;
        mem_45[51]=8'h55;
        mem_45[52]=8'h5c;
        mem_45[53]=8'h5f;
        mem_45[54]=8'h5a;
        mem_45[55]=8'h59;
        mem_45[56]=8'h48;
        mem_45[57]=8'h4b;
        mem_45[58]=8'h4e;
        mem_45[59]=8'h4d;
        mem_45[60]=8'h44;
        mem_45[61]=8'h47;
        mem_45[62]=8'h42;
        mem_45[63]=8'h41;
        mem_45[64]=8'hc0;
        mem_45[65]=8'hc3;
        mem_45[66]=8'hc6;
        mem_45[67]=8'hc5;
        mem_45[68]=8'hcc;
        mem_45[69]=8'hcf;
        mem_45[70]=8'hca;
        mem_45[71]=8'hc9;
        mem_45[72]=8'hd8;
        mem_45[73]=8'hdb;
        mem_45[74]=8'hde;
        mem_45[75]=8'hdd;
        mem_45[76]=8'hd4;
        mem_45[77]=8'hd7;
        mem_45[78]=8'hd2;
        mem_45[79]=8'hd1;
        mem_45[80]=8'hf0;
        mem_45[81]=8'hf3;
        mem_45[82]=8'hf6;
        mem_45[83]=8'hf5;
        mem_45[84]=8'hfc;
        mem_45[85]=8'hff;
        mem_45[86]=8'hfa;
        mem_45[87]=8'hf9;
        mem_45[88]=8'he8;
        mem_45[89]=8'heb;
        mem_45[90]=8'hee;
        mem_45[91]=8'hed;
        mem_45[92]=8'he4;
        mem_45[93]=8'he7;
        mem_45[94]=8'he2;
        mem_45[95]=8'he1;
        mem_45[96]=8'ha0;
        mem_45[97]=8'ha3;
        mem_45[98]=8'ha6;
        mem_45[99]=8'ha5;
        mem_45[100]=8'hac;
        mem_45[101]=8'haf;
        mem_45[102]=8'haa;
        mem_45[103]=8'ha9;
        mem_45[104]=8'hb8;
        mem_45[105]=8'hbb;
        mem_45[106]=8'hbe;
        mem_45[107]=8'hbd;
        mem_45[108]=8'hb4;
        mem_45[109]=8'hb7;
        mem_45[110]=8'hb2;
        mem_45[111]=8'hb1;
        mem_45[112]=8'h90;
        mem_45[113]=8'h93;
        mem_45[114]=8'h96;
        mem_45[115]=8'h95;
        mem_45[116]=8'h9c;
        mem_45[117]=8'h9f;
        mem_45[118]=8'h9a;
        mem_45[119]=8'h99;
        mem_45[120]=8'h88;
        mem_45[121]=8'h8b;
        mem_45[122]=8'h8e;
        mem_45[123]=8'h8d;
        mem_45[124]=8'h84;
        mem_45[125]=8'h87;
        mem_45[126]=8'h82;
        mem_45[127]=8'h81;
        mem_45[128]=8'h9b;
        mem_45[129]=8'h98;
        mem_45[130]=8'h9d;
        mem_45[131]=8'h9e;
        mem_45[132]=8'h97;
        mem_45[133]=8'h94;
        mem_45[134]=8'h91;
        mem_45[135]=8'h92;
        mem_45[136]=8'h83;
        mem_45[137]=8'h80;
        mem_45[138]=8'h85;
        mem_45[139]=8'h86;
        mem_45[140]=8'h8f;
        mem_45[141]=8'h8c;
        mem_45[142]=8'h89;
        mem_45[143]=8'h8a;
        mem_45[144]=8'hab;
        mem_45[145]=8'ha8;
        mem_45[146]=8'had;
        mem_45[147]=8'hae;
        mem_45[148]=8'ha7;
        mem_45[149]=8'ha4;
        mem_45[150]=8'ha1;
        mem_45[151]=8'ha2;
        mem_45[152]=8'hb3;
        mem_45[153]=8'hb0;
        mem_45[154]=8'hb5;
        mem_45[155]=8'hb6;
        mem_45[156]=8'hbf;
        mem_45[157]=8'hbc;
        mem_45[158]=8'hb9;
        mem_45[159]=8'hba;
        mem_45[160]=8'hfb;
        mem_45[161]=8'hf8;
        mem_45[162]=8'hfd;
        mem_45[163]=8'hfe;
        mem_45[164]=8'hf7;
        mem_45[165]=8'hf4;
        mem_45[166]=8'hf1;
        mem_45[167]=8'hf2;
        mem_45[168]=8'he3;
        mem_45[169]=8'he0;
        mem_45[170]=8'he5;
        mem_45[171]=8'he6;
        mem_45[172]=8'hef;
        mem_45[173]=8'hec;
        mem_45[174]=8'he9;
        mem_45[175]=8'hea;
        mem_45[176]=8'hcb;
        mem_45[177]=8'hc8;
        mem_45[178]=8'hcd;
        mem_45[179]=8'hce;
        mem_45[180]=8'hc7;
        mem_45[181]=8'hc4;
        mem_45[182]=8'hc1;
        mem_45[183]=8'hc2;
        mem_45[184]=8'hd3;
        mem_45[185]=8'hd0;
        mem_45[186]=8'hd5;
        mem_45[187]=8'hd6;
        mem_45[188]=8'hdf;
        mem_45[189]=8'hdc;
        mem_45[190]=8'hd9;
        mem_45[191]=8'hda;
        mem_45[192]=8'h5b;
        mem_45[193]=8'h58;
        mem_45[194]=8'h5d;
        mem_45[195]=8'h5e;
        mem_45[196]=8'h57;
        mem_45[197]=8'h54;
        mem_45[198]=8'h51;
        mem_45[199]=8'h52;
        mem_45[200]=8'h43;
        mem_45[201]=8'h40;
        mem_45[202]=8'h45;
        mem_45[203]=8'h46;
        mem_45[204]=8'h4f;
        mem_45[205]=8'h4c;
        mem_45[206]=8'h49;
        mem_45[207]=8'h4a;
        mem_45[208]=8'h6b;
        mem_45[209]=8'h68;
        mem_45[210]=8'h6d;
        mem_45[211]=8'h6e;
        mem_45[212]=8'h67;
        mem_45[213]=8'h64;
        mem_45[214]=8'h61;
        mem_45[215]=8'h62;
        mem_45[216]=8'h73;
        mem_45[217]=8'h70;
        mem_45[218]=8'h75;
        mem_45[219]=8'h76;
        mem_45[220]=8'h7f;
        mem_45[221]=8'h7c;
        mem_45[222]=8'h79;
        mem_45[223]=8'h7a;
        mem_45[224]=8'h3b;
        mem_45[225]=8'h38;
        mem_45[226]=8'h3d;
        mem_45[227]=8'h3e;
        mem_45[228]=8'h37;
        mem_45[229]=8'h34;
        mem_45[230]=8'h31;
        mem_45[231]=8'h32;
        mem_45[232]=8'h23;
        mem_45[233]=8'h20;
        mem_45[234]=8'h25;
        mem_45[235]=8'h26;
        mem_45[236]=8'h2f;
        mem_45[237]=8'h2c;
        mem_45[238]=8'h29;
        mem_45[239]=8'h2a;
        mem_45[240]=8'hb;
        mem_45[241]=8'h8;
        mem_45[242]=8'hd;
        mem_45[243]=8'he;
        mem_45[244]=8'h7;
        mem_45[245]=8'h4;
        mem_45[246]=8'h1;
        mem_45[247]=8'h2;
        mem_45[248]=8'h13;
        mem_45[249]=8'h10;
        mem_45[250]=8'h15;
        mem_45[251]=8'h16;
        mem_45[252]=8'h1f;
        mem_45[253]=8'h1c;
        mem_45[254]=8'h19;
        mem_45[255]=8'h1a;
    end

    initial begin
        mem_46[0]=8'h0;
        mem_46[1]=8'h2;
        mem_46[2]=8'h4;
        mem_46[3]=8'h6;
        mem_46[4]=8'h8;
        mem_46[5]=8'ha;
        mem_46[6]=8'hc;
        mem_46[7]=8'he;
        mem_46[8]=8'h10;
        mem_46[9]=8'h12;
        mem_46[10]=8'h14;
        mem_46[11]=8'h16;
        mem_46[12]=8'h18;
        mem_46[13]=8'h1a;
        mem_46[14]=8'h1c;
        mem_46[15]=8'h1e;
        mem_46[16]=8'h20;
        mem_46[17]=8'h22;
        mem_46[18]=8'h24;
        mem_46[19]=8'h26;
        mem_46[20]=8'h28;
        mem_46[21]=8'h2a;
        mem_46[22]=8'h2c;
        mem_46[23]=8'h2e;
        mem_46[24]=8'h30;
        mem_46[25]=8'h32;
        mem_46[26]=8'h34;
        mem_46[27]=8'h36;
        mem_46[28]=8'h38;
        mem_46[29]=8'h3a;
        mem_46[30]=8'h3c;
        mem_46[31]=8'h3e;
        mem_46[32]=8'h40;
        mem_46[33]=8'h42;
        mem_46[34]=8'h44;
        mem_46[35]=8'h46;
        mem_46[36]=8'h48;
        mem_46[37]=8'h4a;
        mem_46[38]=8'h4c;
        mem_46[39]=8'h4e;
        mem_46[40]=8'h50;
        mem_46[41]=8'h52;
        mem_46[42]=8'h54;
        mem_46[43]=8'h56;
        mem_46[44]=8'h58;
        mem_46[45]=8'h5a;
        mem_46[46]=8'h5c;
        mem_46[47]=8'h5e;
        mem_46[48]=8'h60;
        mem_46[49]=8'h62;
        mem_46[50]=8'h64;
        mem_46[51]=8'h66;
        mem_46[52]=8'h68;
        mem_46[53]=8'h6a;
        mem_46[54]=8'h6c;
        mem_46[55]=8'h6e;
        mem_46[56]=8'h70;
        mem_46[57]=8'h72;
        mem_46[58]=8'h74;
        mem_46[59]=8'h76;
        mem_46[60]=8'h78;
        mem_46[61]=8'h7a;
        mem_46[62]=8'h7c;
        mem_46[63]=8'h7e;
        mem_46[64]=8'h80;
        mem_46[65]=8'h82;
        mem_46[66]=8'h84;
        mem_46[67]=8'h86;
        mem_46[68]=8'h88;
        mem_46[69]=8'h8a;
        mem_46[70]=8'h8c;
        mem_46[71]=8'h8e;
        mem_46[72]=8'h90;
        mem_46[73]=8'h92;
        mem_46[74]=8'h94;
        mem_46[75]=8'h96;
        mem_46[76]=8'h98;
        mem_46[77]=8'h9a;
        mem_46[78]=8'h9c;
        mem_46[79]=8'h9e;
        mem_46[80]=8'ha0;
        mem_46[81]=8'ha2;
        mem_46[82]=8'ha4;
        mem_46[83]=8'ha6;
        mem_46[84]=8'ha8;
        mem_46[85]=8'haa;
        mem_46[86]=8'hac;
        mem_46[87]=8'hae;
        mem_46[88]=8'hb0;
        mem_46[89]=8'hb2;
        mem_46[90]=8'hb4;
        mem_46[91]=8'hb6;
        mem_46[92]=8'hb8;
        mem_46[93]=8'hba;
        mem_46[94]=8'hbc;
        mem_46[95]=8'hbe;
        mem_46[96]=8'hc0;
        mem_46[97]=8'hc2;
        mem_46[98]=8'hc4;
        mem_46[99]=8'hc6;
        mem_46[100]=8'hc8;
        mem_46[101]=8'hca;
        mem_46[102]=8'hcc;
        mem_46[103]=8'hce;
        mem_46[104]=8'hd0;
        mem_46[105]=8'hd2;
        mem_46[106]=8'hd4;
        mem_46[107]=8'hd6;
        mem_46[108]=8'hd8;
        mem_46[109]=8'hda;
        mem_46[110]=8'hdc;
        mem_46[111]=8'hde;
        mem_46[112]=8'he0;
        mem_46[113]=8'he2;
        mem_46[114]=8'he4;
        mem_46[115]=8'he6;
        mem_46[116]=8'he8;
        mem_46[117]=8'hea;
        mem_46[118]=8'hec;
        mem_46[119]=8'hee;
        mem_46[120]=8'hf0;
        mem_46[121]=8'hf2;
        mem_46[122]=8'hf4;
        mem_46[123]=8'hf6;
        mem_46[124]=8'hf8;
        mem_46[125]=8'hfa;
        mem_46[126]=8'hfc;
        mem_46[127]=8'hfe;
        mem_46[128]=8'h1b;
        mem_46[129]=8'h19;
        mem_46[130]=8'h1f;
        mem_46[131]=8'h1d;
        mem_46[132]=8'h13;
        mem_46[133]=8'h11;
        mem_46[134]=8'h17;
        mem_46[135]=8'h15;
        mem_46[136]=8'hb;
        mem_46[137]=8'h9;
        mem_46[138]=8'hf;
        mem_46[139]=8'hd;
        mem_46[140]=8'h3;
        mem_46[141]=8'h1;
        mem_46[142]=8'h7;
        mem_46[143]=8'h5;
        mem_46[144]=8'h3b;
        mem_46[145]=8'h39;
        mem_46[146]=8'h3f;
        mem_46[147]=8'h3d;
        mem_46[148]=8'h33;
        mem_46[149]=8'h31;
        mem_46[150]=8'h37;
        mem_46[151]=8'h35;
        mem_46[152]=8'h2b;
        mem_46[153]=8'h29;
        mem_46[154]=8'h2f;
        mem_46[155]=8'h2d;
        mem_46[156]=8'h23;
        mem_46[157]=8'h21;
        mem_46[158]=8'h27;
        mem_46[159]=8'h25;
        mem_46[160]=8'h5b;
        mem_46[161]=8'h59;
        mem_46[162]=8'h5f;
        mem_46[163]=8'h5d;
        mem_46[164]=8'h53;
        mem_46[165]=8'h51;
        mem_46[166]=8'h57;
        mem_46[167]=8'h55;
        mem_46[168]=8'h4b;
        mem_46[169]=8'h49;
        mem_46[170]=8'h4f;
        mem_46[171]=8'h4d;
        mem_46[172]=8'h43;
        mem_46[173]=8'h41;
        mem_46[174]=8'h47;
        mem_46[175]=8'h45;
        mem_46[176]=8'h7b;
        mem_46[177]=8'h79;
        mem_46[178]=8'h7f;
        mem_46[179]=8'h7d;
        mem_46[180]=8'h73;
        mem_46[181]=8'h71;
        mem_46[182]=8'h77;
        mem_46[183]=8'h75;
        mem_46[184]=8'h6b;
        mem_46[185]=8'h69;
        mem_46[186]=8'h6f;
        mem_46[187]=8'h6d;
        mem_46[188]=8'h63;
        mem_46[189]=8'h61;
        mem_46[190]=8'h67;
        mem_46[191]=8'h65;
        mem_46[192]=8'h9b;
        mem_46[193]=8'h99;
        mem_46[194]=8'h9f;
        mem_46[195]=8'h9d;
        mem_46[196]=8'h93;
        mem_46[197]=8'h91;
        mem_46[198]=8'h97;
        mem_46[199]=8'h95;
        mem_46[200]=8'h8b;
        mem_46[201]=8'h89;
        mem_46[202]=8'h8f;
        mem_46[203]=8'h8d;
        mem_46[204]=8'h83;
        mem_46[205]=8'h81;
        mem_46[206]=8'h87;
        mem_46[207]=8'h85;
        mem_46[208]=8'hbb;
        mem_46[209]=8'hb9;
        mem_46[210]=8'hbf;
        mem_46[211]=8'hbd;
        mem_46[212]=8'hb3;
        mem_46[213]=8'hb1;
        mem_46[214]=8'hb7;
        mem_46[215]=8'hb5;
        mem_46[216]=8'hab;
        mem_46[217]=8'ha9;
        mem_46[218]=8'haf;
        mem_46[219]=8'had;
        mem_46[220]=8'ha3;
        mem_46[221]=8'ha1;
        mem_46[222]=8'ha7;
        mem_46[223]=8'ha5;
        mem_46[224]=8'hdb;
        mem_46[225]=8'hd9;
        mem_46[226]=8'hdf;
        mem_46[227]=8'hdd;
        mem_46[228]=8'hd3;
        mem_46[229]=8'hd1;
        mem_46[230]=8'hd7;
        mem_46[231]=8'hd5;
        mem_46[232]=8'hcb;
        mem_46[233]=8'hc9;
        mem_46[234]=8'hcf;
        mem_46[235]=8'hcd;
        mem_46[236]=8'hc3;
        mem_46[237]=8'hc1;
        mem_46[238]=8'hc7;
        mem_46[239]=8'hc5;
        mem_46[240]=8'hfb;
        mem_46[241]=8'hf9;
        mem_46[242]=8'hff;
        mem_46[243]=8'hfd;
        mem_46[244]=8'hf3;
        mem_46[245]=8'hf1;
        mem_46[246]=8'hf7;
        mem_46[247]=8'hf5;
        mem_46[248]=8'heb;
        mem_46[249]=8'he9;
        mem_46[250]=8'hef;
        mem_46[251]=8'hed;
        mem_46[252]=8'he3;
        mem_46[253]=8'he1;
        mem_46[254]=8'he7;
        mem_46[255]=8'he5;
    end

    initial begin
        mem_47[0]=8'h0;
        mem_47[1]=8'h3;
        mem_47[2]=8'h6;
        mem_47[3]=8'h5;
        mem_47[4]=8'hc;
        mem_47[5]=8'hf;
        mem_47[6]=8'ha;
        mem_47[7]=8'h9;
        mem_47[8]=8'h18;
        mem_47[9]=8'h1b;
        mem_47[10]=8'h1e;
        mem_47[11]=8'h1d;
        mem_47[12]=8'h14;
        mem_47[13]=8'h17;
        mem_47[14]=8'h12;
        mem_47[15]=8'h11;
        mem_47[16]=8'h30;
        mem_47[17]=8'h33;
        mem_47[18]=8'h36;
        mem_47[19]=8'h35;
        mem_47[20]=8'h3c;
        mem_47[21]=8'h3f;
        mem_47[22]=8'h3a;
        mem_47[23]=8'h39;
        mem_47[24]=8'h28;
        mem_47[25]=8'h2b;
        mem_47[26]=8'h2e;
        mem_47[27]=8'h2d;
        mem_47[28]=8'h24;
        mem_47[29]=8'h27;
        mem_47[30]=8'h22;
        mem_47[31]=8'h21;
        mem_47[32]=8'h60;
        mem_47[33]=8'h63;
        mem_47[34]=8'h66;
        mem_47[35]=8'h65;
        mem_47[36]=8'h6c;
        mem_47[37]=8'h6f;
        mem_47[38]=8'h6a;
        mem_47[39]=8'h69;
        mem_47[40]=8'h78;
        mem_47[41]=8'h7b;
        mem_47[42]=8'h7e;
        mem_47[43]=8'h7d;
        mem_47[44]=8'h74;
        mem_47[45]=8'h77;
        mem_47[46]=8'h72;
        mem_47[47]=8'h71;
        mem_47[48]=8'h50;
        mem_47[49]=8'h53;
        mem_47[50]=8'h56;
        mem_47[51]=8'h55;
        mem_47[52]=8'h5c;
        mem_47[53]=8'h5f;
        mem_47[54]=8'h5a;
        mem_47[55]=8'h59;
        mem_47[56]=8'h48;
        mem_47[57]=8'h4b;
        mem_47[58]=8'h4e;
        mem_47[59]=8'h4d;
        mem_47[60]=8'h44;
        mem_47[61]=8'h47;
        mem_47[62]=8'h42;
        mem_47[63]=8'h41;
        mem_47[64]=8'hc0;
        mem_47[65]=8'hc3;
        mem_47[66]=8'hc6;
        mem_47[67]=8'hc5;
        mem_47[68]=8'hcc;
        mem_47[69]=8'hcf;
        mem_47[70]=8'hca;
        mem_47[71]=8'hc9;
        mem_47[72]=8'hd8;
        mem_47[73]=8'hdb;
        mem_47[74]=8'hde;
        mem_47[75]=8'hdd;
        mem_47[76]=8'hd4;
        mem_47[77]=8'hd7;
        mem_47[78]=8'hd2;
        mem_47[79]=8'hd1;
        mem_47[80]=8'hf0;
        mem_47[81]=8'hf3;
        mem_47[82]=8'hf6;
        mem_47[83]=8'hf5;
        mem_47[84]=8'hfc;
        mem_47[85]=8'hff;
        mem_47[86]=8'hfa;
        mem_47[87]=8'hf9;
        mem_47[88]=8'he8;
        mem_47[89]=8'heb;
        mem_47[90]=8'hee;
        mem_47[91]=8'hed;
        mem_47[92]=8'he4;
        mem_47[93]=8'he7;
        mem_47[94]=8'he2;
        mem_47[95]=8'he1;
        mem_47[96]=8'ha0;
        mem_47[97]=8'ha3;
        mem_47[98]=8'ha6;
        mem_47[99]=8'ha5;
        mem_47[100]=8'hac;
        mem_47[101]=8'haf;
        mem_47[102]=8'haa;
        mem_47[103]=8'ha9;
        mem_47[104]=8'hb8;
        mem_47[105]=8'hbb;
        mem_47[106]=8'hbe;
        mem_47[107]=8'hbd;
        mem_47[108]=8'hb4;
        mem_47[109]=8'hb7;
        mem_47[110]=8'hb2;
        mem_47[111]=8'hb1;
        mem_47[112]=8'h90;
        mem_47[113]=8'h93;
        mem_47[114]=8'h96;
        mem_47[115]=8'h95;
        mem_47[116]=8'h9c;
        mem_47[117]=8'h9f;
        mem_47[118]=8'h9a;
        mem_47[119]=8'h99;
        mem_47[120]=8'h88;
        mem_47[121]=8'h8b;
        mem_47[122]=8'h8e;
        mem_47[123]=8'h8d;
        mem_47[124]=8'h84;
        mem_47[125]=8'h87;
        mem_47[126]=8'h82;
        mem_47[127]=8'h81;
        mem_47[128]=8'h9b;
        mem_47[129]=8'h98;
        mem_47[130]=8'h9d;
        mem_47[131]=8'h9e;
        mem_47[132]=8'h97;
        mem_47[133]=8'h94;
        mem_47[134]=8'h91;
        mem_47[135]=8'h92;
        mem_47[136]=8'h83;
        mem_47[137]=8'h80;
        mem_47[138]=8'h85;
        mem_47[139]=8'h86;
        mem_47[140]=8'h8f;
        mem_47[141]=8'h8c;
        mem_47[142]=8'h89;
        mem_47[143]=8'h8a;
        mem_47[144]=8'hab;
        mem_47[145]=8'ha8;
        mem_47[146]=8'had;
        mem_47[147]=8'hae;
        mem_47[148]=8'ha7;
        mem_47[149]=8'ha4;
        mem_47[150]=8'ha1;
        mem_47[151]=8'ha2;
        mem_47[152]=8'hb3;
        mem_47[153]=8'hb0;
        mem_47[154]=8'hb5;
        mem_47[155]=8'hb6;
        mem_47[156]=8'hbf;
        mem_47[157]=8'hbc;
        mem_47[158]=8'hb9;
        mem_47[159]=8'hba;
        mem_47[160]=8'hfb;
        mem_47[161]=8'hf8;
        mem_47[162]=8'hfd;
        mem_47[163]=8'hfe;
        mem_47[164]=8'hf7;
        mem_47[165]=8'hf4;
        mem_47[166]=8'hf1;
        mem_47[167]=8'hf2;
        mem_47[168]=8'he3;
        mem_47[169]=8'he0;
        mem_47[170]=8'he5;
        mem_47[171]=8'he6;
        mem_47[172]=8'hef;
        mem_47[173]=8'hec;
        mem_47[174]=8'he9;
        mem_47[175]=8'hea;
        mem_47[176]=8'hcb;
        mem_47[177]=8'hc8;
        mem_47[178]=8'hcd;
        mem_47[179]=8'hce;
        mem_47[180]=8'hc7;
        mem_47[181]=8'hc4;
        mem_47[182]=8'hc1;
        mem_47[183]=8'hc2;
        mem_47[184]=8'hd3;
        mem_47[185]=8'hd0;
        mem_47[186]=8'hd5;
        mem_47[187]=8'hd6;
        mem_47[188]=8'hdf;
        mem_47[189]=8'hdc;
        mem_47[190]=8'hd9;
        mem_47[191]=8'hda;
        mem_47[192]=8'h5b;
        mem_47[193]=8'h58;
        mem_47[194]=8'h5d;
        mem_47[195]=8'h5e;
        mem_47[196]=8'h57;
        mem_47[197]=8'h54;
        mem_47[198]=8'h51;
        mem_47[199]=8'h52;
        mem_47[200]=8'h43;
        mem_47[201]=8'h40;
        mem_47[202]=8'h45;
        mem_47[203]=8'h46;
        mem_47[204]=8'h4f;
        mem_47[205]=8'h4c;
        mem_47[206]=8'h49;
        mem_47[207]=8'h4a;
        mem_47[208]=8'h6b;
        mem_47[209]=8'h68;
        mem_47[210]=8'h6d;
        mem_47[211]=8'h6e;
        mem_47[212]=8'h67;
        mem_47[213]=8'h64;
        mem_47[214]=8'h61;
        mem_47[215]=8'h62;
        mem_47[216]=8'h73;
        mem_47[217]=8'h70;
        mem_47[218]=8'h75;
        mem_47[219]=8'h76;
        mem_47[220]=8'h7f;
        mem_47[221]=8'h7c;
        mem_47[222]=8'h79;
        mem_47[223]=8'h7a;
        mem_47[224]=8'h3b;
        mem_47[225]=8'h38;
        mem_47[226]=8'h3d;
        mem_47[227]=8'h3e;
        mem_47[228]=8'h37;
        mem_47[229]=8'h34;
        mem_47[230]=8'h31;
        mem_47[231]=8'h32;
        mem_47[232]=8'h23;
        mem_47[233]=8'h20;
        mem_47[234]=8'h25;
        mem_47[235]=8'h26;
        mem_47[236]=8'h2f;
        mem_47[237]=8'h2c;
        mem_47[238]=8'h29;
        mem_47[239]=8'h2a;
        mem_47[240]=8'hb;
        mem_47[241]=8'h8;
        mem_47[242]=8'hd;
        mem_47[243]=8'he;
        mem_47[244]=8'h7;
        mem_47[245]=8'h4;
        mem_47[246]=8'h1;
        mem_47[247]=8'h2;
        mem_47[248]=8'h13;
        mem_47[249]=8'h10;
        mem_47[250]=8'h15;
        mem_47[251]=8'h16;
        mem_47[252]=8'h1f;
        mem_47[253]=8'h1c;
        mem_47[254]=8'h19;
        mem_47[255]=8'h1a;
    end

    initial begin
        mem_48[0]=8'h0;
        mem_48[1]=8'h2;
        mem_48[2]=8'h4;
        mem_48[3]=8'h6;
        mem_48[4]=8'h8;
        mem_48[5]=8'ha;
        mem_48[6]=8'hc;
        mem_48[7]=8'he;
        mem_48[8]=8'h10;
        mem_48[9]=8'h12;
        mem_48[10]=8'h14;
        mem_48[11]=8'h16;
        mem_48[12]=8'h18;
        mem_48[13]=8'h1a;
        mem_48[14]=8'h1c;
        mem_48[15]=8'h1e;
        mem_48[16]=8'h20;
        mem_48[17]=8'h22;
        mem_48[18]=8'h24;
        mem_48[19]=8'h26;
        mem_48[20]=8'h28;
        mem_48[21]=8'h2a;
        mem_48[22]=8'h2c;
        mem_48[23]=8'h2e;
        mem_48[24]=8'h30;
        mem_48[25]=8'h32;
        mem_48[26]=8'h34;
        mem_48[27]=8'h36;
        mem_48[28]=8'h38;
        mem_48[29]=8'h3a;
        mem_48[30]=8'h3c;
        mem_48[31]=8'h3e;
        mem_48[32]=8'h40;
        mem_48[33]=8'h42;
        mem_48[34]=8'h44;
        mem_48[35]=8'h46;
        mem_48[36]=8'h48;
        mem_48[37]=8'h4a;
        mem_48[38]=8'h4c;
        mem_48[39]=8'h4e;
        mem_48[40]=8'h50;
        mem_48[41]=8'h52;
        mem_48[42]=8'h54;
        mem_48[43]=8'h56;
        mem_48[44]=8'h58;
        mem_48[45]=8'h5a;
        mem_48[46]=8'h5c;
        mem_48[47]=8'h5e;
        mem_48[48]=8'h60;
        mem_48[49]=8'h62;
        mem_48[50]=8'h64;
        mem_48[51]=8'h66;
        mem_48[52]=8'h68;
        mem_48[53]=8'h6a;
        mem_48[54]=8'h6c;
        mem_48[55]=8'h6e;
        mem_48[56]=8'h70;
        mem_48[57]=8'h72;
        mem_48[58]=8'h74;
        mem_48[59]=8'h76;
        mem_48[60]=8'h78;
        mem_48[61]=8'h7a;
        mem_48[62]=8'h7c;
        mem_48[63]=8'h7e;
        mem_48[64]=8'h80;
        mem_48[65]=8'h82;
        mem_48[66]=8'h84;
        mem_48[67]=8'h86;
        mem_48[68]=8'h88;
        mem_48[69]=8'h8a;
        mem_48[70]=8'h8c;
        mem_48[71]=8'h8e;
        mem_48[72]=8'h90;
        mem_48[73]=8'h92;
        mem_48[74]=8'h94;
        mem_48[75]=8'h96;
        mem_48[76]=8'h98;
        mem_48[77]=8'h9a;
        mem_48[78]=8'h9c;
        mem_48[79]=8'h9e;
        mem_48[80]=8'ha0;
        mem_48[81]=8'ha2;
        mem_48[82]=8'ha4;
        mem_48[83]=8'ha6;
        mem_48[84]=8'ha8;
        mem_48[85]=8'haa;
        mem_48[86]=8'hac;
        mem_48[87]=8'hae;
        mem_48[88]=8'hb0;
        mem_48[89]=8'hb2;
        mem_48[90]=8'hb4;
        mem_48[91]=8'hb6;
        mem_48[92]=8'hb8;
        mem_48[93]=8'hba;
        mem_48[94]=8'hbc;
        mem_48[95]=8'hbe;
        mem_48[96]=8'hc0;
        mem_48[97]=8'hc2;
        mem_48[98]=8'hc4;
        mem_48[99]=8'hc6;
        mem_48[100]=8'hc8;
        mem_48[101]=8'hca;
        mem_48[102]=8'hcc;
        mem_48[103]=8'hce;
        mem_48[104]=8'hd0;
        mem_48[105]=8'hd2;
        mem_48[106]=8'hd4;
        mem_48[107]=8'hd6;
        mem_48[108]=8'hd8;
        mem_48[109]=8'hda;
        mem_48[110]=8'hdc;
        mem_48[111]=8'hde;
        mem_48[112]=8'he0;
        mem_48[113]=8'he2;
        mem_48[114]=8'he4;
        mem_48[115]=8'he6;
        mem_48[116]=8'he8;
        mem_48[117]=8'hea;
        mem_48[118]=8'hec;
        mem_48[119]=8'hee;
        mem_48[120]=8'hf0;
        mem_48[121]=8'hf2;
        mem_48[122]=8'hf4;
        mem_48[123]=8'hf6;
        mem_48[124]=8'hf8;
        mem_48[125]=8'hfa;
        mem_48[126]=8'hfc;
        mem_48[127]=8'hfe;
        mem_48[128]=8'h1b;
        mem_48[129]=8'h19;
        mem_48[130]=8'h1f;
        mem_48[131]=8'h1d;
        mem_48[132]=8'h13;
        mem_48[133]=8'h11;
        mem_48[134]=8'h17;
        mem_48[135]=8'h15;
        mem_48[136]=8'hb;
        mem_48[137]=8'h9;
        mem_48[138]=8'hf;
        mem_48[139]=8'hd;
        mem_48[140]=8'h3;
        mem_48[141]=8'h1;
        mem_48[142]=8'h7;
        mem_48[143]=8'h5;
        mem_48[144]=8'h3b;
        mem_48[145]=8'h39;
        mem_48[146]=8'h3f;
        mem_48[147]=8'h3d;
        mem_48[148]=8'h33;
        mem_48[149]=8'h31;
        mem_48[150]=8'h37;
        mem_48[151]=8'h35;
        mem_48[152]=8'h2b;
        mem_48[153]=8'h29;
        mem_48[154]=8'h2f;
        mem_48[155]=8'h2d;
        mem_48[156]=8'h23;
        mem_48[157]=8'h21;
        mem_48[158]=8'h27;
        mem_48[159]=8'h25;
        mem_48[160]=8'h5b;
        mem_48[161]=8'h59;
        mem_48[162]=8'h5f;
        mem_48[163]=8'h5d;
        mem_48[164]=8'h53;
        mem_48[165]=8'h51;
        mem_48[166]=8'h57;
        mem_48[167]=8'h55;
        mem_48[168]=8'h4b;
        mem_48[169]=8'h49;
        mem_48[170]=8'h4f;
        mem_48[171]=8'h4d;
        mem_48[172]=8'h43;
        mem_48[173]=8'h41;
        mem_48[174]=8'h47;
        mem_48[175]=8'h45;
        mem_48[176]=8'h7b;
        mem_48[177]=8'h79;
        mem_48[178]=8'h7f;
        mem_48[179]=8'h7d;
        mem_48[180]=8'h73;
        mem_48[181]=8'h71;
        mem_48[182]=8'h77;
        mem_48[183]=8'h75;
        mem_48[184]=8'h6b;
        mem_48[185]=8'h69;
        mem_48[186]=8'h6f;
        mem_48[187]=8'h6d;
        mem_48[188]=8'h63;
        mem_48[189]=8'h61;
        mem_48[190]=8'h67;
        mem_48[191]=8'h65;
        mem_48[192]=8'h9b;
        mem_48[193]=8'h99;
        mem_48[194]=8'h9f;
        mem_48[195]=8'h9d;
        mem_48[196]=8'h93;
        mem_48[197]=8'h91;
        mem_48[198]=8'h97;
        mem_48[199]=8'h95;
        mem_48[200]=8'h8b;
        mem_48[201]=8'h89;
        mem_48[202]=8'h8f;
        mem_48[203]=8'h8d;
        mem_48[204]=8'h83;
        mem_48[205]=8'h81;
        mem_48[206]=8'h87;
        mem_48[207]=8'h85;
        mem_48[208]=8'hbb;
        mem_48[209]=8'hb9;
        mem_48[210]=8'hbf;
        mem_48[211]=8'hbd;
        mem_48[212]=8'hb3;
        mem_48[213]=8'hb1;
        mem_48[214]=8'hb7;
        mem_48[215]=8'hb5;
        mem_48[216]=8'hab;
        mem_48[217]=8'ha9;
        mem_48[218]=8'haf;
        mem_48[219]=8'had;
        mem_48[220]=8'ha3;
        mem_48[221]=8'ha1;
        mem_48[222]=8'ha7;
        mem_48[223]=8'ha5;
        mem_48[224]=8'hdb;
        mem_48[225]=8'hd9;
        mem_48[226]=8'hdf;
        mem_48[227]=8'hdd;
        mem_48[228]=8'hd3;
        mem_48[229]=8'hd1;
        mem_48[230]=8'hd7;
        mem_48[231]=8'hd5;
        mem_48[232]=8'hcb;
        mem_48[233]=8'hc9;
        mem_48[234]=8'hcf;
        mem_48[235]=8'hcd;
        mem_48[236]=8'hc3;
        mem_48[237]=8'hc1;
        mem_48[238]=8'hc7;
        mem_48[239]=8'hc5;
        mem_48[240]=8'hfb;
        mem_48[241]=8'hf9;
        mem_48[242]=8'hff;
        mem_48[243]=8'hfd;
        mem_48[244]=8'hf3;
        mem_48[245]=8'hf1;
        mem_48[246]=8'hf7;
        mem_48[247]=8'hf5;
        mem_48[248]=8'heb;
        mem_48[249]=8'he9;
        mem_48[250]=8'hef;
        mem_48[251]=8'hed;
        mem_48[252]=8'he3;
        mem_48[253]=8'he1;
        mem_48[254]=8'he7;
        mem_48[255]=8'he5;
    end

    initial begin
        mem_49[0]=8'h0;
        mem_49[1]=8'h3;
        mem_49[2]=8'h6;
        mem_49[3]=8'h5;
        mem_49[4]=8'hc;
        mem_49[5]=8'hf;
        mem_49[6]=8'ha;
        mem_49[7]=8'h9;
        mem_49[8]=8'h18;
        mem_49[9]=8'h1b;
        mem_49[10]=8'h1e;
        mem_49[11]=8'h1d;
        mem_49[12]=8'h14;
        mem_49[13]=8'h17;
        mem_49[14]=8'h12;
        mem_49[15]=8'h11;
        mem_49[16]=8'h30;
        mem_49[17]=8'h33;
        mem_49[18]=8'h36;
        mem_49[19]=8'h35;
        mem_49[20]=8'h3c;
        mem_49[21]=8'h3f;
        mem_49[22]=8'h3a;
        mem_49[23]=8'h39;
        mem_49[24]=8'h28;
        mem_49[25]=8'h2b;
        mem_49[26]=8'h2e;
        mem_49[27]=8'h2d;
        mem_49[28]=8'h24;
        mem_49[29]=8'h27;
        mem_49[30]=8'h22;
        mem_49[31]=8'h21;
        mem_49[32]=8'h60;
        mem_49[33]=8'h63;
        mem_49[34]=8'h66;
        mem_49[35]=8'h65;
        mem_49[36]=8'h6c;
        mem_49[37]=8'h6f;
        mem_49[38]=8'h6a;
        mem_49[39]=8'h69;
        mem_49[40]=8'h78;
        mem_49[41]=8'h7b;
        mem_49[42]=8'h7e;
        mem_49[43]=8'h7d;
        mem_49[44]=8'h74;
        mem_49[45]=8'h77;
        mem_49[46]=8'h72;
        mem_49[47]=8'h71;
        mem_49[48]=8'h50;
        mem_49[49]=8'h53;
        mem_49[50]=8'h56;
        mem_49[51]=8'h55;
        mem_49[52]=8'h5c;
        mem_49[53]=8'h5f;
        mem_49[54]=8'h5a;
        mem_49[55]=8'h59;
        mem_49[56]=8'h48;
        mem_49[57]=8'h4b;
        mem_49[58]=8'h4e;
        mem_49[59]=8'h4d;
        mem_49[60]=8'h44;
        mem_49[61]=8'h47;
        mem_49[62]=8'h42;
        mem_49[63]=8'h41;
        mem_49[64]=8'hc0;
        mem_49[65]=8'hc3;
        mem_49[66]=8'hc6;
        mem_49[67]=8'hc5;
        mem_49[68]=8'hcc;
        mem_49[69]=8'hcf;
        mem_49[70]=8'hca;
        mem_49[71]=8'hc9;
        mem_49[72]=8'hd8;
        mem_49[73]=8'hdb;
        mem_49[74]=8'hde;
        mem_49[75]=8'hdd;
        mem_49[76]=8'hd4;
        mem_49[77]=8'hd7;
        mem_49[78]=8'hd2;
        mem_49[79]=8'hd1;
        mem_49[80]=8'hf0;
        mem_49[81]=8'hf3;
        mem_49[82]=8'hf6;
        mem_49[83]=8'hf5;
        mem_49[84]=8'hfc;
        mem_49[85]=8'hff;
        mem_49[86]=8'hfa;
        mem_49[87]=8'hf9;
        mem_49[88]=8'he8;
        mem_49[89]=8'heb;
        mem_49[90]=8'hee;
        mem_49[91]=8'hed;
        mem_49[92]=8'he4;
        mem_49[93]=8'he7;
        mem_49[94]=8'he2;
        mem_49[95]=8'he1;
        mem_49[96]=8'ha0;
        mem_49[97]=8'ha3;
        mem_49[98]=8'ha6;
        mem_49[99]=8'ha5;
        mem_49[100]=8'hac;
        mem_49[101]=8'haf;
        mem_49[102]=8'haa;
        mem_49[103]=8'ha9;
        mem_49[104]=8'hb8;
        mem_49[105]=8'hbb;
        mem_49[106]=8'hbe;
        mem_49[107]=8'hbd;
        mem_49[108]=8'hb4;
        mem_49[109]=8'hb7;
        mem_49[110]=8'hb2;
        mem_49[111]=8'hb1;
        mem_49[112]=8'h90;
        mem_49[113]=8'h93;
        mem_49[114]=8'h96;
        mem_49[115]=8'h95;
        mem_49[116]=8'h9c;
        mem_49[117]=8'h9f;
        mem_49[118]=8'h9a;
        mem_49[119]=8'h99;
        mem_49[120]=8'h88;
        mem_49[121]=8'h8b;
        mem_49[122]=8'h8e;
        mem_49[123]=8'h8d;
        mem_49[124]=8'h84;
        mem_49[125]=8'h87;
        mem_49[126]=8'h82;
        mem_49[127]=8'h81;
        mem_49[128]=8'h9b;
        mem_49[129]=8'h98;
        mem_49[130]=8'h9d;
        mem_49[131]=8'h9e;
        mem_49[132]=8'h97;
        mem_49[133]=8'h94;
        mem_49[134]=8'h91;
        mem_49[135]=8'h92;
        mem_49[136]=8'h83;
        mem_49[137]=8'h80;
        mem_49[138]=8'h85;
        mem_49[139]=8'h86;
        mem_49[140]=8'h8f;
        mem_49[141]=8'h8c;
        mem_49[142]=8'h89;
        mem_49[143]=8'h8a;
        mem_49[144]=8'hab;
        mem_49[145]=8'ha8;
        mem_49[146]=8'had;
        mem_49[147]=8'hae;
        mem_49[148]=8'ha7;
        mem_49[149]=8'ha4;
        mem_49[150]=8'ha1;
        mem_49[151]=8'ha2;
        mem_49[152]=8'hb3;
        mem_49[153]=8'hb0;
        mem_49[154]=8'hb5;
        mem_49[155]=8'hb6;
        mem_49[156]=8'hbf;
        mem_49[157]=8'hbc;
        mem_49[158]=8'hb9;
        mem_49[159]=8'hba;
        mem_49[160]=8'hfb;
        mem_49[161]=8'hf8;
        mem_49[162]=8'hfd;
        mem_49[163]=8'hfe;
        mem_49[164]=8'hf7;
        mem_49[165]=8'hf4;
        mem_49[166]=8'hf1;
        mem_49[167]=8'hf2;
        mem_49[168]=8'he3;
        mem_49[169]=8'he0;
        mem_49[170]=8'he5;
        mem_49[171]=8'he6;
        mem_49[172]=8'hef;
        mem_49[173]=8'hec;
        mem_49[174]=8'he9;
        mem_49[175]=8'hea;
        mem_49[176]=8'hcb;
        mem_49[177]=8'hc8;
        mem_49[178]=8'hcd;
        mem_49[179]=8'hce;
        mem_49[180]=8'hc7;
        mem_49[181]=8'hc4;
        mem_49[182]=8'hc1;
        mem_49[183]=8'hc2;
        mem_49[184]=8'hd3;
        mem_49[185]=8'hd0;
        mem_49[186]=8'hd5;
        mem_49[187]=8'hd6;
        mem_49[188]=8'hdf;
        mem_49[189]=8'hdc;
        mem_49[190]=8'hd9;
        mem_49[191]=8'hda;
        mem_49[192]=8'h5b;
        mem_49[193]=8'h58;
        mem_49[194]=8'h5d;
        mem_49[195]=8'h5e;
        mem_49[196]=8'h57;
        mem_49[197]=8'h54;
        mem_49[198]=8'h51;
        mem_49[199]=8'h52;
        mem_49[200]=8'h43;
        mem_49[201]=8'h40;
        mem_49[202]=8'h45;
        mem_49[203]=8'h46;
        mem_49[204]=8'h4f;
        mem_49[205]=8'h4c;
        mem_49[206]=8'h49;
        mem_49[207]=8'h4a;
        mem_49[208]=8'h6b;
        mem_49[209]=8'h68;
        mem_49[210]=8'h6d;
        mem_49[211]=8'h6e;
        mem_49[212]=8'h67;
        mem_49[213]=8'h64;
        mem_49[214]=8'h61;
        mem_49[215]=8'h62;
        mem_49[216]=8'h73;
        mem_49[217]=8'h70;
        mem_49[218]=8'h75;
        mem_49[219]=8'h76;
        mem_49[220]=8'h7f;
        mem_49[221]=8'h7c;
        mem_49[222]=8'h79;
        mem_49[223]=8'h7a;
        mem_49[224]=8'h3b;
        mem_49[225]=8'h38;
        mem_49[226]=8'h3d;
        mem_49[227]=8'h3e;
        mem_49[228]=8'h37;
        mem_49[229]=8'h34;
        mem_49[230]=8'h31;
        mem_49[231]=8'h32;
        mem_49[232]=8'h23;
        mem_49[233]=8'h20;
        mem_49[234]=8'h25;
        mem_49[235]=8'h26;
        mem_49[236]=8'h2f;
        mem_49[237]=8'h2c;
        mem_49[238]=8'h29;
        mem_49[239]=8'h2a;
        mem_49[240]=8'hb;
        mem_49[241]=8'h8;
        mem_49[242]=8'hd;
        mem_49[243]=8'he;
        mem_49[244]=8'h7;
        mem_49[245]=8'h4;
        mem_49[246]=8'h1;
        mem_49[247]=8'h2;
        mem_49[248]=8'h13;
        mem_49[249]=8'h10;
        mem_49[250]=8'h15;
        mem_49[251]=8'h16;
        mem_49[252]=8'h1f;
        mem_49[253]=8'h1c;
        mem_49[254]=8'h19;
        mem_49[255]=8'h1a;
    end

    initial begin
        mem_50[0]=8'h0;
        mem_50[1]=8'h2;
        mem_50[2]=8'h4;
        mem_50[3]=8'h6;
        mem_50[4]=8'h8;
        mem_50[5]=8'ha;
        mem_50[6]=8'hc;
        mem_50[7]=8'he;
        mem_50[8]=8'h10;
        mem_50[9]=8'h12;
        mem_50[10]=8'h14;
        mem_50[11]=8'h16;
        mem_50[12]=8'h18;
        mem_50[13]=8'h1a;
        mem_50[14]=8'h1c;
        mem_50[15]=8'h1e;
        mem_50[16]=8'h20;
        mem_50[17]=8'h22;
        mem_50[18]=8'h24;
        mem_50[19]=8'h26;
        mem_50[20]=8'h28;
        mem_50[21]=8'h2a;
        mem_50[22]=8'h2c;
        mem_50[23]=8'h2e;
        mem_50[24]=8'h30;
        mem_50[25]=8'h32;
        mem_50[26]=8'h34;
        mem_50[27]=8'h36;
        mem_50[28]=8'h38;
        mem_50[29]=8'h3a;
        mem_50[30]=8'h3c;
        mem_50[31]=8'h3e;
        mem_50[32]=8'h40;
        mem_50[33]=8'h42;
        mem_50[34]=8'h44;
        mem_50[35]=8'h46;
        mem_50[36]=8'h48;
        mem_50[37]=8'h4a;
        mem_50[38]=8'h4c;
        mem_50[39]=8'h4e;
        mem_50[40]=8'h50;
        mem_50[41]=8'h52;
        mem_50[42]=8'h54;
        mem_50[43]=8'h56;
        mem_50[44]=8'h58;
        mem_50[45]=8'h5a;
        mem_50[46]=8'h5c;
        mem_50[47]=8'h5e;
        mem_50[48]=8'h60;
        mem_50[49]=8'h62;
        mem_50[50]=8'h64;
        mem_50[51]=8'h66;
        mem_50[52]=8'h68;
        mem_50[53]=8'h6a;
        mem_50[54]=8'h6c;
        mem_50[55]=8'h6e;
        mem_50[56]=8'h70;
        mem_50[57]=8'h72;
        mem_50[58]=8'h74;
        mem_50[59]=8'h76;
        mem_50[60]=8'h78;
        mem_50[61]=8'h7a;
        mem_50[62]=8'h7c;
        mem_50[63]=8'h7e;
        mem_50[64]=8'h80;
        mem_50[65]=8'h82;
        mem_50[66]=8'h84;
        mem_50[67]=8'h86;
        mem_50[68]=8'h88;
        mem_50[69]=8'h8a;
        mem_50[70]=8'h8c;
        mem_50[71]=8'h8e;
        mem_50[72]=8'h90;
        mem_50[73]=8'h92;
        mem_50[74]=8'h94;
        mem_50[75]=8'h96;
        mem_50[76]=8'h98;
        mem_50[77]=8'h9a;
        mem_50[78]=8'h9c;
        mem_50[79]=8'h9e;
        mem_50[80]=8'ha0;
        mem_50[81]=8'ha2;
        mem_50[82]=8'ha4;
        mem_50[83]=8'ha6;
        mem_50[84]=8'ha8;
        mem_50[85]=8'haa;
        mem_50[86]=8'hac;
        mem_50[87]=8'hae;
        mem_50[88]=8'hb0;
        mem_50[89]=8'hb2;
        mem_50[90]=8'hb4;
        mem_50[91]=8'hb6;
        mem_50[92]=8'hb8;
        mem_50[93]=8'hba;
        mem_50[94]=8'hbc;
        mem_50[95]=8'hbe;
        mem_50[96]=8'hc0;
        mem_50[97]=8'hc2;
        mem_50[98]=8'hc4;
        mem_50[99]=8'hc6;
        mem_50[100]=8'hc8;
        mem_50[101]=8'hca;
        mem_50[102]=8'hcc;
        mem_50[103]=8'hce;
        mem_50[104]=8'hd0;
        mem_50[105]=8'hd2;
        mem_50[106]=8'hd4;
        mem_50[107]=8'hd6;
        mem_50[108]=8'hd8;
        mem_50[109]=8'hda;
        mem_50[110]=8'hdc;
        mem_50[111]=8'hde;
        mem_50[112]=8'he0;
        mem_50[113]=8'he2;
        mem_50[114]=8'he4;
        mem_50[115]=8'he6;
        mem_50[116]=8'he8;
        mem_50[117]=8'hea;
        mem_50[118]=8'hec;
        mem_50[119]=8'hee;
        mem_50[120]=8'hf0;
        mem_50[121]=8'hf2;
        mem_50[122]=8'hf4;
        mem_50[123]=8'hf6;
        mem_50[124]=8'hf8;
        mem_50[125]=8'hfa;
        mem_50[126]=8'hfc;
        mem_50[127]=8'hfe;
        mem_50[128]=8'h1b;
        mem_50[129]=8'h19;
        mem_50[130]=8'h1f;
        mem_50[131]=8'h1d;
        mem_50[132]=8'h13;
        mem_50[133]=8'h11;
        mem_50[134]=8'h17;
        mem_50[135]=8'h15;
        mem_50[136]=8'hb;
        mem_50[137]=8'h9;
        mem_50[138]=8'hf;
        mem_50[139]=8'hd;
        mem_50[140]=8'h3;
        mem_50[141]=8'h1;
        mem_50[142]=8'h7;
        mem_50[143]=8'h5;
        mem_50[144]=8'h3b;
        mem_50[145]=8'h39;
        mem_50[146]=8'h3f;
        mem_50[147]=8'h3d;
        mem_50[148]=8'h33;
        mem_50[149]=8'h31;
        mem_50[150]=8'h37;
        mem_50[151]=8'h35;
        mem_50[152]=8'h2b;
        mem_50[153]=8'h29;
        mem_50[154]=8'h2f;
        mem_50[155]=8'h2d;
        mem_50[156]=8'h23;
        mem_50[157]=8'h21;
        mem_50[158]=8'h27;
        mem_50[159]=8'h25;
        mem_50[160]=8'h5b;
        mem_50[161]=8'h59;
        mem_50[162]=8'h5f;
        mem_50[163]=8'h5d;
        mem_50[164]=8'h53;
        mem_50[165]=8'h51;
        mem_50[166]=8'h57;
        mem_50[167]=8'h55;
        mem_50[168]=8'h4b;
        mem_50[169]=8'h49;
        mem_50[170]=8'h4f;
        mem_50[171]=8'h4d;
        mem_50[172]=8'h43;
        mem_50[173]=8'h41;
        mem_50[174]=8'h47;
        mem_50[175]=8'h45;
        mem_50[176]=8'h7b;
        mem_50[177]=8'h79;
        mem_50[178]=8'h7f;
        mem_50[179]=8'h7d;
        mem_50[180]=8'h73;
        mem_50[181]=8'h71;
        mem_50[182]=8'h77;
        mem_50[183]=8'h75;
        mem_50[184]=8'h6b;
        mem_50[185]=8'h69;
        mem_50[186]=8'h6f;
        mem_50[187]=8'h6d;
        mem_50[188]=8'h63;
        mem_50[189]=8'h61;
        mem_50[190]=8'h67;
        mem_50[191]=8'h65;
        mem_50[192]=8'h9b;
        mem_50[193]=8'h99;
        mem_50[194]=8'h9f;
        mem_50[195]=8'h9d;
        mem_50[196]=8'h93;
        mem_50[197]=8'h91;
        mem_50[198]=8'h97;
        mem_50[199]=8'h95;
        mem_50[200]=8'h8b;
        mem_50[201]=8'h89;
        mem_50[202]=8'h8f;
        mem_50[203]=8'h8d;
        mem_50[204]=8'h83;
        mem_50[205]=8'h81;
        mem_50[206]=8'h87;
        mem_50[207]=8'h85;
        mem_50[208]=8'hbb;
        mem_50[209]=8'hb9;
        mem_50[210]=8'hbf;
        mem_50[211]=8'hbd;
        mem_50[212]=8'hb3;
        mem_50[213]=8'hb1;
        mem_50[214]=8'hb7;
        mem_50[215]=8'hb5;
        mem_50[216]=8'hab;
        mem_50[217]=8'ha9;
        mem_50[218]=8'haf;
        mem_50[219]=8'had;
        mem_50[220]=8'ha3;
        mem_50[221]=8'ha1;
        mem_50[222]=8'ha7;
        mem_50[223]=8'ha5;
        mem_50[224]=8'hdb;
        mem_50[225]=8'hd9;
        mem_50[226]=8'hdf;
        mem_50[227]=8'hdd;
        mem_50[228]=8'hd3;
        mem_50[229]=8'hd1;
        mem_50[230]=8'hd7;
        mem_50[231]=8'hd5;
        mem_50[232]=8'hcb;
        mem_50[233]=8'hc9;
        mem_50[234]=8'hcf;
        mem_50[235]=8'hcd;
        mem_50[236]=8'hc3;
        mem_50[237]=8'hc1;
        mem_50[238]=8'hc7;
        mem_50[239]=8'hc5;
        mem_50[240]=8'hfb;
        mem_50[241]=8'hf9;
        mem_50[242]=8'hff;
        mem_50[243]=8'hfd;
        mem_50[244]=8'hf3;
        mem_50[245]=8'hf1;
        mem_50[246]=8'hf7;
        mem_50[247]=8'hf5;
        mem_50[248]=8'heb;
        mem_50[249]=8'he9;
        mem_50[250]=8'hef;
        mem_50[251]=8'hed;
        mem_50[252]=8'he3;
        mem_50[253]=8'he1;
        mem_50[254]=8'he7;
        mem_50[255]=8'he5;
    end

    initial begin
        mem_51[0]=8'h0;
        mem_51[1]=8'h3;
        mem_51[2]=8'h6;
        mem_51[3]=8'h5;
        mem_51[4]=8'hc;
        mem_51[5]=8'hf;
        mem_51[6]=8'ha;
        mem_51[7]=8'h9;
        mem_51[8]=8'h18;
        mem_51[9]=8'h1b;
        mem_51[10]=8'h1e;
        mem_51[11]=8'h1d;
        mem_51[12]=8'h14;
        mem_51[13]=8'h17;
        mem_51[14]=8'h12;
        mem_51[15]=8'h11;
        mem_51[16]=8'h30;
        mem_51[17]=8'h33;
        mem_51[18]=8'h36;
        mem_51[19]=8'h35;
        mem_51[20]=8'h3c;
        mem_51[21]=8'h3f;
        mem_51[22]=8'h3a;
        mem_51[23]=8'h39;
        mem_51[24]=8'h28;
        mem_51[25]=8'h2b;
        mem_51[26]=8'h2e;
        mem_51[27]=8'h2d;
        mem_51[28]=8'h24;
        mem_51[29]=8'h27;
        mem_51[30]=8'h22;
        mem_51[31]=8'h21;
        mem_51[32]=8'h60;
        mem_51[33]=8'h63;
        mem_51[34]=8'h66;
        mem_51[35]=8'h65;
        mem_51[36]=8'h6c;
        mem_51[37]=8'h6f;
        mem_51[38]=8'h6a;
        mem_51[39]=8'h69;
        mem_51[40]=8'h78;
        mem_51[41]=8'h7b;
        mem_51[42]=8'h7e;
        mem_51[43]=8'h7d;
        mem_51[44]=8'h74;
        mem_51[45]=8'h77;
        mem_51[46]=8'h72;
        mem_51[47]=8'h71;
        mem_51[48]=8'h50;
        mem_51[49]=8'h53;
        mem_51[50]=8'h56;
        mem_51[51]=8'h55;
        mem_51[52]=8'h5c;
        mem_51[53]=8'h5f;
        mem_51[54]=8'h5a;
        mem_51[55]=8'h59;
        mem_51[56]=8'h48;
        mem_51[57]=8'h4b;
        mem_51[58]=8'h4e;
        mem_51[59]=8'h4d;
        mem_51[60]=8'h44;
        mem_51[61]=8'h47;
        mem_51[62]=8'h42;
        mem_51[63]=8'h41;
        mem_51[64]=8'hc0;
        mem_51[65]=8'hc3;
        mem_51[66]=8'hc6;
        mem_51[67]=8'hc5;
        mem_51[68]=8'hcc;
        mem_51[69]=8'hcf;
        mem_51[70]=8'hca;
        mem_51[71]=8'hc9;
        mem_51[72]=8'hd8;
        mem_51[73]=8'hdb;
        mem_51[74]=8'hde;
        mem_51[75]=8'hdd;
        mem_51[76]=8'hd4;
        mem_51[77]=8'hd7;
        mem_51[78]=8'hd2;
        mem_51[79]=8'hd1;
        mem_51[80]=8'hf0;
        mem_51[81]=8'hf3;
        mem_51[82]=8'hf6;
        mem_51[83]=8'hf5;
        mem_51[84]=8'hfc;
        mem_51[85]=8'hff;
        mem_51[86]=8'hfa;
        mem_51[87]=8'hf9;
        mem_51[88]=8'he8;
        mem_51[89]=8'heb;
        mem_51[90]=8'hee;
        mem_51[91]=8'hed;
        mem_51[92]=8'he4;
        mem_51[93]=8'he7;
        mem_51[94]=8'he2;
        mem_51[95]=8'he1;
        mem_51[96]=8'ha0;
        mem_51[97]=8'ha3;
        mem_51[98]=8'ha6;
        mem_51[99]=8'ha5;
        mem_51[100]=8'hac;
        mem_51[101]=8'haf;
        mem_51[102]=8'haa;
        mem_51[103]=8'ha9;
        mem_51[104]=8'hb8;
        mem_51[105]=8'hbb;
        mem_51[106]=8'hbe;
        mem_51[107]=8'hbd;
        mem_51[108]=8'hb4;
        mem_51[109]=8'hb7;
        mem_51[110]=8'hb2;
        mem_51[111]=8'hb1;
        mem_51[112]=8'h90;
        mem_51[113]=8'h93;
        mem_51[114]=8'h96;
        mem_51[115]=8'h95;
        mem_51[116]=8'h9c;
        mem_51[117]=8'h9f;
        mem_51[118]=8'h9a;
        mem_51[119]=8'h99;
        mem_51[120]=8'h88;
        mem_51[121]=8'h8b;
        mem_51[122]=8'h8e;
        mem_51[123]=8'h8d;
        mem_51[124]=8'h84;
        mem_51[125]=8'h87;
        mem_51[126]=8'h82;
        mem_51[127]=8'h81;
        mem_51[128]=8'h9b;
        mem_51[129]=8'h98;
        mem_51[130]=8'h9d;
        mem_51[131]=8'h9e;
        mem_51[132]=8'h97;
        mem_51[133]=8'h94;
        mem_51[134]=8'h91;
        mem_51[135]=8'h92;
        mem_51[136]=8'h83;
        mem_51[137]=8'h80;
        mem_51[138]=8'h85;
        mem_51[139]=8'h86;
        mem_51[140]=8'h8f;
        mem_51[141]=8'h8c;
        mem_51[142]=8'h89;
        mem_51[143]=8'h8a;
        mem_51[144]=8'hab;
        mem_51[145]=8'ha8;
        mem_51[146]=8'had;
        mem_51[147]=8'hae;
        mem_51[148]=8'ha7;
        mem_51[149]=8'ha4;
        mem_51[150]=8'ha1;
        mem_51[151]=8'ha2;
        mem_51[152]=8'hb3;
        mem_51[153]=8'hb0;
        mem_51[154]=8'hb5;
        mem_51[155]=8'hb6;
        mem_51[156]=8'hbf;
        mem_51[157]=8'hbc;
        mem_51[158]=8'hb9;
        mem_51[159]=8'hba;
        mem_51[160]=8'hfb;
        mem_51[161]=8'hf8;
        mem_51[162]=8'hfd;
        mem_51[163]=8'hfe;
        mem_51[164]=8'hf7;
        mem_51[165]=8'hf4;
        mem_51[166]=8'hf1;
        mem_51[167]=8'hf2;
        mem_51[168]=8'he3;
        mem_51[169]=8'he0;
        mem_51[170]=8'he5;
        mem_51[171]=8'he6;
        mem_51[172]=8'hef;
        mem_51[173]=8'hec;
        mem_51[174]=8'he9;
        mem_51[175]=8'hea;
        mem_51[176]=8'hcb;
        mem_51[177]=8'hc8;
        mem_51[178]=8'hcd;
        mem_51[179]=8'hce;
        mem_51[180]=8'hc7;
        mem_51[181]=8'hc4;
        mem_51[182]=8'hc1;
        mem_51[183]=8'hc2;
        mem_51[184]=8'hd3;
        mem_51[185]=8'hd0;
        mem_51[186]=8'hd5;
        mem_51[187]=8'hd6;
        mem_51[188]=8'hdf;
        mem_51[189]=8'hdc;
        mem_51[190]=8'hd9;
        mem_51[191]=8'hda;
        mem_51[192]=8'h5b;
        mem_51[193]=8'h58;
        mem_51[194]=8'h5d;
        mem_51[195]=8'h5e;
        mem_51[196]=8'h57;
        mem_51[197]=8'h54;
        mem_51[198]=8'h51;
        mem_51[199]=8'h52;
        mem_51[200]=8'h43;
        mem_51[201]=8'h40;
        mem_51[202]=8'h45;
        mem_51[203]=8'h46;
        mem_51[204]=8'h4f;
        mem_51[205]=8'h4c;
        mem_51[206]=8'h49;
        mem_51[207]=8'h4a;
        mem_51[208]=8'h6b;
        mem_51[209]=8'h68;
        mem_51[210]=8'h6d;
        mem_51[211]=8'h6e;
        mem_51[212]=8'h67;
        mem_51[213]=8'h64;
        mem_51[214]=8'h61;
        mem_51[215]=8'h62;
        mem_51[216]=8'h73;
        mem_51[217]=8'h70;
        mem_51[218]=8'h75;
        mem_51[219]=8'h76;
        mem_51[220]=8'h7f;
        mem_51[221]=8'h7c;
        mem_51[222]=8'h79;
        mem_51[223]=8'h7a;
        mem_51[224]=8'h3b;
        mem_51[225]=8'h38;
        mem_51[226]=8'h3d;
        mem_51[227]=8'h3e;
        mem_51[228]=8'h37;
        mem_51[229]=8'h34;
        mem_51[230]=8'h31;
        mem_51[231]=8'h32;
        mem_51[232]=8'h23;
        mem_51[233]=8'h20;
        mem_51[234]=8'h25;
        mem_51[235]=8'h26;
        mem_51[236]=8'h2f;
        mem_51[237]=8'h2c;
        mem_51[238]=8'h29;
        mem_51[239]=8'h2a;
        mem_51[240]=8'hb;
        mem_51[241]=8'h8;
        mem_51[242]=8'hd;
        mem_51[243]=8'he;
        mem_51[244]=8'h7;
        mem_51[245]=8'h4;
        mem_51[246]=8'h1;
        mem_51[247]=8'h2;
        mem_51[248]=8'h13;
        mem_51[249]=8'h10;
        mem_51[250]=8'h15;
        mem_51[251]=8'h16;
        mem_51[252]=8'h1f;
        mem_51[253]=8'h1c;
        mem_51[254]=8'h19;
        mem_51[255]=8'h1a;
    end

    initial begin
        mem_52[0]=8'h0;
        mem_52[1]=8'h2;
        mem_52[2]=8'h4;
        mem_52[3]=8'h6;
        mem_52[4]=8'h8;
        mem_52[5]=8'ha;
        mem_52[6]=8'hc;
        mem_52[7]=8'he;
        mem_52[8]=8'h10;
        mem_52[9]=8'h12;
        mem_52[10]=8'h14;
        mem_52[11]=8'h16;
        mem_52[12]=8'h18;
        mem_52[13]=8'h1a;
        mem_52[14]=8'h1c;
        mem_52[15]=8'h1e;
        mem_52[16]=8'h20;
        mem_52[17]=8'h22;
        mem_52[18]=8'h24;
        mem_52[19]=8'h26;
        mem_52[20]=8'h28;
        mem_52[21]=8'h2a;
        mem_52[22]=8'h2c;
        mem_52[23]=8'h2e;
        mem_52[24]=8'h30;
        mem_52[25]=8'h32;
        mem_52[26]=8'h34;
        mem_52[27]=8'h36;
        mem_52[28]=8'h38;
        mem_52[29]=8'h3a;
        mem_52[30]=8'h3c;
        mem_52[31]=8'h3e;
        mem_52[32]=8'h40;
        mem_52[33]=8'h42;
        mem_52[34]=8'h44;
        mem_52[35]=8'h46;
        mem_52[36]=8'h48;
        mem_52[37]=8'h4a;
        mem_52[38]=8'h4c;
        mem_52[39]=8'h4e;
        mem_52[40]=8'h50;
        mem_52[41]=8'h52;
        mem_52[42]=8'h54;
        mem_52[43]=8'h56;
        mem_52[44]=8'h58;
        mem_52[45]=8'h5a;
        mem_52[46]=8'h5c;
        mem_52[47]=8'h5e;
        mem_52[48]=8'h60;
        mem_52[49]=8'h62;
        mem_52[50]=8'h64;
        mem_52[51]=8'h66;
        mem_52[52]=8'h68;
        mem_52[53]=8'h6a;
        mem_52[54]=8'h6c;
        mem_52[55]=8'h6e;
        mem_52[56]=8'h70;
        mem_52[57]=8'h72;
        mem_52[58]=8'h74;
        mem_52[59]=8'h76;
        mem_52[60]=8'h78;
        mem_52[61]=8'h7a;
        mem_52[62]=8'h7c;
        mem_52[63]=8'h7e;
        mem_52[64]=8'h80;
        mem_52[65]=8'h82;
        mem_52[66]=8'h84;
        mem_52[67]=8'h86;
        mem_52[68]=8'h88;
        mem_52[69]=8'h8a;
        mem_52[70]=8'h8c;
        mem_52[71]=8'h8e;
        mem_52[72]=8'h90;
        mem_52[73]=8'h92;
        mem_52[74]=8'h94;
        mem_52[75]=8'h96;
        mem_52[76]=8'h98;
        mem_52[77]=8'h9a;
        mem_52[78]=8'h9c;
        mem_52[79]=8'h9e;
        mem_52[80]=8'ha0;
        mem_52[81]=8'ha2;
        mem_52[82]=8'ha4;
        mem_52[83]=8'ha6;
        mem_52[84]=8'ha8;
        mem_52[85]=8'haa;
        mem_52[86]=8'hac;
        mem_52[87]=8'hae;
        mem_52[88]=8'hb0;
        mem_52[89]=8'hb2;
        mem_52[90]=8'hb4;
        mem_52[91]=8'hb6;
        mem_52[92]=8'hb8;
        mem_52[93]=8'hba;
        mem_52[94]=8'hbc;
        mem_52[95]=8'hbe;
        mem_52[96]=8'hc0;
        mem_52[97]=8'hc2;
        mem_52[98]=8'hc4;
        mem_52[99]=8'hc6;
        mem_52[100]=8'hc8;
        mem_52[101]=8'hca;
        mem_52[102]=8'hcc;
        mem_52[103]=8'hce;
        mem_52[104]=8'hd0;
        mem_52[105]=8'hd2;
        mem_52[106]=8'hd4;
        mem_52[107]=8'hd6;
        mem_52[108]=8'hd8;
        mem_52[109]=8'hda;
        mem_52[110]=8'hdc;
        mem_52[111]=8'hde;
        mem_52[112]=8'he0;
        mem_52[113]=8'he2;
        mem_52[114]=8'he4;
        mem_52[115]=8'he6;
        mem_52[116]=8'he8;
        mem_52[117]=8'hea;
        mem_52[118]=8'hec;
        mem_52[119]=8'hee;
        mem_52[120]=8'hf0;
        mem_52[121]=8'hf2;
        mem_52[122]=8'hf4;
        mem_52[123]=8'hf6;
        mem_52[124]=8'hf8;
        mem_52[125]=8'hfa;
        mem_52[126]=8'hfc;
        mem_52[127]=8'hfe;
        mem_52[128]=8'h1b;
        mem_52[129]=8'h19;
        mem_52[130]=8'h1f;
        mem_52[131]=8'h1d;
        mem_52[132]=8'h13;
        mem_52[133]=8'h11;
        mem_52[134]=8'h17;
        mem_52[135]=8'h15;
        mem_52[136]=8'hb;
        mem_52[137]=8'h9;
        mem_52[138]=8'hf;
        mem_52[139]=8'hd;
        mem_52[140]=8'h3;
        mem_52[141]=8'h1;
        mem_52[142]=8'h7;
        mem_52[143]=8'h5;
        mem_52[144]=8'h3b;
        mem_52[145]=8'h39;
        mem_52[146]=8'h3f;
        mem_52[147]=8'h3d;
        mem_52[148]=8'h33;
        mem_52[149]=8'h31;
        mem_52[150]=8'h37;
        mem_52[151]=8'h35;
        mem_52[152]=8'h2b;
        mem_52[153]=8'h29;
        mem_52[154]=8'h2f;
        mem_52[155]=8'h2d;
        mem_52[156]=8'h23;
        mem_52[157]=8'h21;
        mem_52[158]=8'h27;
        mem_52[159]=8'h25;
        mem_52[160]=8'h5b;
        mem_52[161]=8'h59;
        mem_52[162]=8'h5f;
        mem_52[163]=8'h5d;
        mem_52[164]=8'h53;
        mem_52[165]=8'h51;
        mem_52[166]=8'h57;
        mem_52[167]=8'h55;
        mem_52[168]=8'h4b;
        mem_52[169]=8'h49;
        mem_52[170]=8'h4f;
        mem_52[171]=8'h4d;
        mem_52[172]=8'h43;
        mem_52[173]=8'h41;
        mem_52[174]=8'h47;
        mem_52[175]=8'h45;
        mem_52[176]=8'h7b;
        mem_52[177]=8'h79;
        mem_52[178]=8'h7f;
        mem_52[179]=8'h7d;
        mem_52[180]=8'h73;
        mem_52[181]=8'h71;
        mem_52[182]=8'h77;
        mem_52[183]=8'h75;
        mem_52[184]=8'h6b;
        mem_52[185]=8'h69;
        mem_52[186]=8'h6f;
        mem_52[187]=8'h6d;
        mem_52[188]=8'h63;
        mem_52[189]=8'h61;
        mem_52[190]=8'h67;
        mem_52[191]=8'h65;
        mem_52[192]=8'h9b;
        mem_52[193]=8'h99;
        mem_52[194]=8'h9f;
        mem_52[195]=8'h9d;
        mem_52[196]=8'h93;
        mem_52[197]=8'h91;
        mem_52[198]=8'h97;
        mem_52[199]=8'h95;
        mem_52[200]=8'h8b;
        mem_52[201]=8'h89;
        mem_52[202]=8'h8f;
        mem_52[203]=8'h8d;
        mem_52[204]=8'h83;
        mem_52[205]=8'h81;
        mem_52[206]=8'h87;
        mem_52[207]=8'h85;
        mem_52[208]=8'hbb;
        mem_52[209]=8'hb9;
        mem_52[210]=8'hbf;
        mem_52[211]=8'hbd;
        mem_52[212]=8'hb3;
        mem_52[213]=8'hb1;
        mem_52[214]=8'hb7;
        mem_52[215]=8'hb5;
        mem_52[216]=8'hab;
        mem_52[217]=8'ha9;
        mem_52[218]=8'haf;
        mem_52[219]=8'had;
        mem_52[220]=8'ha3;
        mem_52[221]=8'ha1;
        mem_52[222]=8'ha7;
        mem_52[223]=8'ha5;
        mem_52[224]=8'hdb;
        mem_52[225]=8'hd9;
        mem_52[226]=8'hdf;
        mem_52[227]=8'hdd;
        mem_52[228]=8'hd3;
        mem_52[229]=8'hd1;
        mem_52[230]=8'hd7;
        mem_52[231]=8'hd5;
        mem_52[232]=8'hcb;
        mem_52[233]=8'hc9;
        mem_52[234]=8'hcf;
        mem_52[235]=8'hcd;
        mem_52[236]=8'hc3;
        mem_52[237]=8'hc1;
        mem_52[238]=8'hc7;
        mem_52[239]=8'hc5;
        mem_52[240]=8'hfb;
        mem_52[241]=8'hf9;
        mem_52[242]=8'hff;
        mem_52[243]=8'hfd;
        mem_52[244]=8'hf3;
        mem_52[245]=8'hf1;
        mem_52[246]=8'hf7;
        mem_52[247]=8'hf5;
        mem_52[248]=8'heb;
        mem_52[249]=8'he9;
        mem_52[250]=8'hef;
        mem_52[251]=8'hed;
        mem_52[252]=8'he3;
        mem_52[253]=8'he1;
        mem_52[254]=8'he7;
        mem_52[255]=8'he5;
    end

    initial begin
        mem_53[0]=8'h0;
        mem_53[1]=8'h3;
        mem_53[2]=8'h6;
        mem_53[3]=8'h5;
        mem_53[4]=8'hc;
        mem_53[5]=8'hf;
        mem_53[6]=8'ha;
        mem_53[7]=8'h9;
        mem_53[8]=8'h18;
        mem_53[9]=8'h1b;
        mem_53[10]=8'h1e;
        mem_53[11]=8'h1d;
        mem_53[12]=8'h14;
        mem_53[13]=8'h17;
        mem_53[14]=8'h12;
        mem_53[15]=8'h11;
        mem_53[16]=8'h30;
        mem_53[17]=8'h33;
        mem_53[18]=8'h36;
        mem_53[19]=8'h35;
        mem_53[20]=8'h3c;
        mem_53[21]=8'h3f;
        mem_53[22]=8'h3a;
        mem_53[23]=8'h39;
        mem_53[24]=8'h28;
        mem_53[25]=8'h2b;
        mem_53[26]=8'h2e;
        mem_53[27]=8'h2d;
        mem_53[28]=8'h24;
        mem_53[29]=8'h27;
        mem_53[30]=8'h22;
        mem_53[31]=8'h21;
        mem_53[32]=8'h60;
        mem_53[33]=8'h63;
        mem_53[34]=8'h66;
        mem_53[35]=8'h65;
        mem_53[36]=8'h6c;
        mem_53[37]=8'h6f;
        mem_53[38]=8'h6a;
        mem_53[39]=8'h69;
        mem_53[40]=8'h78;
        mem_53[41]=8'h7b;
        mem_53[42]=8'h7e;
        mem_53[43]=8'h7d;
        mem_53[44]=8'h74;
        mem_53[45]=8'h77;
        mem_53[46]=8'h72;
        mem_53[47]=8'h71;
        mem_53[48]=8'h50;
        mem_53[49]=8'h53;
        mem_53[50]=8'h56;
        mem_53[51]=8'h55;
        mem_53[52]=8'h5c;
        mem_53[53]=8'h5f;
        mem_53[54]=8'h5a;
        mem_53[55]=8'h59;
        mem_53[56]=8'h48;
        mem_53[57]=8'h4b;
        mem_53[58]=8'h4e;
        mem_53[59]=8'h4d;
        mem_53[60]=8'h44;
        mem_53[61]=8'h47;
        mem_53[62]=8'h42;
        mem_53[63]=8'h41;
        mem_53[64]=8'hc0;
        mem_53[65]=8'hc3;
        mem_53[66]=8'hc6;
        mem_53[67]=8'hc5;
        mem_53[68]=8'hcc;
        mem_53[69]=8'hcf;
        mem_53[70]=8'hca;
        mem_53[71]=8'hc9;
        mem_53[72]=8'hd8;
        mem_53[73]=8'hdb;
        mem_53[74]=8'hde;
        mem_53[75]=8'hdd;
        mem_53[76]=8'hd4;
        mem_53[77]=8'hd7;
        mem_53[78]=8'hd2;
        mem_53[79]=8'hd1;
        mem_53[80]=8'hf0;
        mem_53[81]=8'hf3;
        mem_53[82]=8'hf6;
        mem_53[83]=8'hf5;
        mem_53[84]=8'hfc;
        mem_53[85]=8'hff;
        mem_53[86]=8'hfa;
        mem_53[87]=8'hf9;
        mem_53[88]=8'he8;
        mem_53[89]=8'heb;
        mem_53[90]=8'hee;
        mem_53[91]=8'hed;
        mem_53[92]=8'he4;
        mem_53[93]=8'he7;
        mem_53[94]=8'he2;
        mem_53[95]=8'he1;
        mem_53[96]=8'ha0;
        mem_53[97]=8'ha3;
        mem_53[98]=8'ha6;
        mem_53[99]=8'ha5;
        mem_53[100]=8'hac;
        mem_53[101]=8'haf;
        mem_53[102]=8'haa;
        mem_53[103]=8'ha9;
        mem_53[104]=8'hb8;
        mem_53[105]=8'hbb;
        mem_53[106]=8'hbe;
        mem_53[107]=8'hbd;
        mem_53[108]=8'hb4;
        mem_53[109]=8'hb7;
        mem_53[110]=8'hb2;
        mem_53[111]=8'hb1;
        mem_53[112]=8'h90;
        mem_53[113]=8'h93;
        mem_53[114]=8'h96;
        mem_53[115]=8'h95;
        mem_53[116]=8'h9c;
        mem_53[117]=8'h9f;
        mem_53[118]=8'h9a;
        mem_53[119]=8'h99;
        mem_53[120]=8'h88;
        mem_53[121]=8'h8b;
        mem_53[122]=8'h8e;
        mem_53[123]=8'h8d;
        mem_53[124]=8'h84;
        mem_53[125]=8'h87;
        mem_53[126]=8'h82;
        mem_53[127]=8'h81;
        mem_53[128]=8'h9b;
        mem_53[129]=8'h98;
        mem_53[130]=8'h9d;
        mem_53[131]=8'h9e;
        mem_53[132]=8'h97;
        mem_53[133]=8'h94;
        mem_53[134]=8'h91;
        mem_53[135]=8'h92;
        mem_53[136]=8'h83;
        mem_53[137]=8'h80;
        mem_53[138]=8'h85;
        mem_53[139]=8'h86;
        mem_53[140]=8'h8f;
        mem_53[141]=8'h8c;
        mem_53[142]=8'h89;
        mem_53[143]=8'h8a;
        mem_53[144]=8'hab;
        mem_53[145]=8'ha8;
        mem_53[146]=8'had;
        mem_53[147]=8'hae;
        mem_53[148]=8'ha7;
        mem_53[149]=8'ha4;
        mem_53[150]=8'ha1;
        mem_53[151]=8'ha2;
        mem_53[152]=8'hb3;
        mem_53[153]=8'hb0;
        mem_53[154]=8'hb5;
        mem_53[155]=8'hb6;
        mem_53[156]=8'hbf;
        mem_53[157]=8'hbc;
        mem_53[158]=8'hb9;
        mem_53[159]=8'hba;
        mem_53[160]=8'hfb;
        mem_53[161]=8'hf8;
        mem_53[162]=8'hfd;
        mem_53[163]=8'hfe;
        mem_53[164]=8'hf7;
        mem_53[165]=8'hf4;
        mem_53[166]=8'hf1;
        mem_53[167]=8'hf2;
        mem_53[168]=8'he3;
        mem_53[169]=8'he0;
        mem_53[170]=8'he5;
        mem_53[171]=8'he6;
        mem_53[172]=8'hef;
        mem_53[173]=8'hec;
        mem_53[174]=8'he9;
        mem_53[175]=8'hea;
        mem_53[176]=8'hcb;
        mem_53[177]=8'hc8;
        mem_53[178]=8'hcd;
        mem_53[179]=8'hce;
        mem_53[180]=8'hc7;
        mem_53[181]=8'hc4;
        mem_53[182]=8'hc1;
        mem_53[183]=8'hc2;
        mem_53[184]=8'hd3;
        mem_53[185]=8'hd0;
        mem_53[186]=8'hd5;
        mem_53[187]=8'hd6;
        mem_53[188]=8'hdf;
        mem_53[189]=8'hdc;
        mem_53[190]=8'hd9;
        mem_53[191]=8'hda;
        mem_53[192]=8'h5b;
        mem_53[193]=8'h58;
        mem_53[194]=8'h5d;
        mem_53[195]=8'h5e;
        mem_53[196]=8'h57;
        mem_53[197]=8'h54;
        mem_53[198]=8'h51;
        mem_53[199]=8'h52;
        mem_53[200]=8'h43;
        mem_53[201]=8'h40;
        mem_53[202]=8'h45;
        mem_53[203]=8'h46;
        mem_53[204]=8'h4f;
        mem_53[205]=8'h4c;
        mem_53[206]=8'h49;
        mem_53[207]=8'h4a;
        mem_53[208]=8'h6b;
        mem_53[209]=8'h68;
        mem_53[210]=8'h6d;
        mem_53[211]=8'h6e;
        mem_53[212]=8'h67;
        mem_53[213]=8'h64;
        mem_53[214]=8'h61;
        mem_53[215]=8'h62;
        mem_53[216]=8'h73;
        mem_53[217]=8'h70;
        mem_53[218]=8'h75;
        mem_53[219]=8'h76;
        mem_53[220]=8'h7f;
        mem_53[221]=8'h7c;
        mem_53[222]=8'h79;
        mem_53[223]=8'h7a;
        mem_53[224]=8'h3b;
        mem_53[225]=8'h38;
        mem_53[226]=8'h3d;
        mem_53[227]=8'h3e;
        mem_53[228]=8'h37;
        mem_53[229]=8'h34;
        mem_53[230]=8'h31;
        mem_53[231]=8'h32;
        mem_53[232]=8'h23;
        mem_53[233]=8'h20;
        mem_53[234]=8'h25;
        mem_53[235]=8'h26;
        mem_53[236]=8'h2f;
        mem_53[237]=8'h2c;
        mem_53[238]=8'h29;
        mem_53[239]=8'h2a;
        mem_53[240]=8'hb;
        mem_53[241]=8'h8;
        mem_53[242]=8'hd;
        mem_53[243]=8'he;
        mem_53[244]=8'h7;
        mem_53[245]=8'h4;
        mem_53[246]=8'h1;
        mem_53[247]=8'h2;
        mem_53[248]=8'h13;
        mem_53[249]=8'h10;
        mem_53[250]=8'h15;
        mem_53[251]=8'h16;
        mem_53[252]=8'h1f;
        mem_53[253]=8'h1c;
        mem_53[254]=8'h19;
        mem_53[255]=8'h1a;
    end

    initial begin
        mem_54[0]=8'h63;
        mem_54[1]=8'h7c;
        mem_54[2]=8'h77;
        mem_54[3]=8'h7b;
        mem_54[4]=8'hf2;
        mem_54[5]=8'h6b;
        mem_54[6]=8'h6f;
        mem_54[7]=8'hc5;
        mem_54[8]=8'h30;
        mem_54[9]=8'h1;
        mem_54[10]=8'h67;
        mem_54[11]=8'h2b;
        mem_54[12]=8'hfe;
        mem_54[13]=8'hd7;
        mem_54[14]=8'hab;
        mem_54[15]=8'h76;
        mem_54[16]=8'hca;
        mem_54[17]=8'h82;
        mem_54[18]=8'hc9;
        mem_54[19]=8'h7d;
        mem_54[20]=8'hfa;
        mem_54[21]=8'h59;
        mem_54[22]=8'h47;
        mem_54[23]=8'hf0;
        mem_54[24]=8'had;
        mem_54[25]=8'hd4;
        mem_54[26]=8'ha2;
        mem_54[27]=8'haf;
        mem_54[28]=8'h9c;
        mem_54[29]=8'ha4;
        mem_54[30]=8'h72;
        mem_54[31]=8'hc0;
        mem_54[32]=8'hb7;
        mem_54[33]=8'hfd;
        mem_54[34]=8'h93;
        mem_54[35]=8'h26;
        mem_54[36]=8'h36;
        mem_54[37]=8'h3f;
        mem_54[38]=8'hf7;
        mem_54[39]=8'hcc;
        mem_54[40]=8'h34;
        mem_54[41]=8'ha5;
        mem_54[42]=8'he5;
        mem_54[43]=8'hf1;
        mem_54[44]=8'h71;
        mem_54[45]=8'hd8;
        mem_54[46]=8'h31;
        mem_54[47]=8'h15;
        mem_54[48]=8'h4;
        mem_54[49]=8'hc7;
        mem_54[50]=8'h23;
        mem_54[51]=8'hc3;
        mem_54[52]=8'h18;
        mem_54[53]=8'h96;
        mem_54[54]=8'h5;
        mem_54[55]=8'h9a;
        mem_54[56]=8'h7;
        mem_54[57]=8'h12;
        mem_54[58]=8'h80;
        mem_54[59]=8'he2;
        mem_54[60]=8'heb;
        mem_54[61]=8'h27;
        mem_54[62]=8'hb2;
        mem_54[63]=8'h75;
        mem_54[64]=8'h9;
        mem_54[65]=8'h83;
        mem_54[66]=8'h2c;
        mem_54[67]=8'h1a;
        mem_54[68]=8'h1b;
        mem_54[69]=8'h6e;
        mem_54[70]=8'h5a;
        mem_54[71]=8'ha0;
        mem_54[72]=8'h52;
        mem_54[73]=8'h3b;
        mem_54[74]=8'hd6;
        mem_54[75]=8'hb3;
        mem_54[76]=8'h29;
        mem_54[77]=8'he3;
        mem_54[78]=8'h2f;
        mem_54[79]=8'h84;
        mem_54[80]=8'h53;
        mem_54[81]=8'hd1;
        mem_54[82]=8'h0;
        mem_54[83]=8'hed;
        mem_54[84]=8'h20;
        mem_54[85]=8'hfc;
        mem_54[86]=8'hb1;
        mem_54[87]=8'h5b;
        mem_54[88]=8'h6a;
        mem_54[89]=8'hcb;
        mem_54[90]=8'hbe;
        mem_54[91]=8'h39;
        mem_54[92]=8'h4a;
        mem_54[93]=8'h4c;
        mem_54[94]=8'h58;
        mem_54[95]=8'hcf;
        mem_54[96]=8'hd0;
        mem_54[97]=8'hef;
        mem_54[98]=8'haa;
        mem_54[99]=8'hfb;
        mem_54[100]=8'h43;
        mem_54[101]=8'h4d;
        mem_54[102]=8'h33;
        mem_54[103]=8'h85;
        mem_54[104]=8'h45;
        mem_54[105]=8'hf9;
        mem_54[106]=8'h2;
        mem_54[107]=8'h7f;
        mem_54[108]=8'h50;
        mem_54[109]=8'h3c;
        mem_54[110]=8'h9f;
        mem_54[111]=8'ha8;
        mem_54[112]=8'h51;
        mem_54[113]=8'ha3;
        mem_54[114]=8'h40;
        mem_54[115]=8'h8f;
        mem_54[116]=8'h92;
        mem_54[117]=8'h9d;
        mem_54[118]=8'h38;
        mem_54[119]=8'hf5;
        mem_54[120]=8'hbc;
        mem_54[121]=8'hb6;
        mem_54[122]=8'hda;
        mem_54[123]=8'h21;
        mem_54[124]=8'h10;
        mem_54[125]=8'hff;
        mem_54[126]=8'hf3;
        mem_54[127]=8'hd2;
        mem_54[128]=8'hcd;
        mem_54[129]=8'hc;
        mem_54[130]=8'h13;
        mem_54[131]=8'hec;
        mem_54[132]=8'h5f;
        mem_54[133]=8'h97;
        mem_54[134]=8'h44;
        mem_54[135]=8'h17;
        mem_54[136]=8'hc4;
        mem_54[137]=8'ha7;
        mem_54[138]=8'h7e;
        mem_54[139]=8'h3d;
        mem_54[140]=8'h64;
        mem_54[141]=8'h5d;
        mem_54[142]=8'h19;
        mem_54[143]=8'h73;
        mem_54[144]=8'h60;
        mem_54[145]=8'h81;
        mem_54[146]=8'h4f;
        mem_54[147]=8'hdc;
        mem_54[148]=8'h22;
        mem_54[149]=8'h2a;
        mem_54[150]=8'h90;
        mem_54[151]=8'h88;
        mem_54[152]=8'h46;
        mem_54[153]=8'hee;
        mem_54[154]=8'hb8;
        mem_54[155]=8'h14;
        mem_54[156]=8'hde;
        mem_54[157]=8'h5e;
        mem_54[158]=8'hb;
        mem_54[159]=8'hdb;
        mem_54[160]=8'he0;
        mem_54[161]=8'h32;
        mem_54[162]=8'h3a;
        mem_54[163]=8'ha;
        mem_54[164]=8'h49;
        mem_54[165]=8'h6;
        mem_54[166]=8'h24;
        mem_54[167]=8'h5c;
        mem_54[168]=8'hc2;
        mem_54[169]=8'hd3;
        mem_54[170]=8'hac;
        mem_54[171]=8'h62;
        mem_54[172]=8'h91;
        mem_54[173]=8'h95;
        mem_54[174]=8'he4;
        mem_54[175]=8'h79;
        mem_54[176]=8'he7;
        mem_54[177]=8'hc8;
        mem_54[178]=8'h37;
        mem_54[179]=8'h6d;
        mem_54[180]=8'h8d;
        mem_54[181]=8'hd5;
        mem_54[182]=8'h4e;
        mem_54[183]=8'ha9;
        mem_54[184]=8'h6c;
        mem_54[185]=8'h56;
        mem_54[186]=8'hf4;
        mem_54[187]=8'hea;
        mem_54[188]=8'h65;
        mem_54[189]=8'h7a;
        mem_54[190]=8'hae;
        mem_54[191]=8'h8;
        mem_54[192]=8'hba;
        mem_54[193]=8'h78;
        mem_54[194]=8'h25;
        mem_54[195]=8'h2e;
        mem_54[196]=8'h1c;
        mem_54[197]=8'ha6;
        mem_54[198]=8'hb4;
        mem_54[199]=8'hc6;
        mem_54[200]=8'he8;
        mem_54[201]=8'hdd;
        mem_54[202]=8'h74;
        mem_54[203]=8'h1f;
        mem_54[204]=8'h4b;
        mem_54[205]=8'hbd;
        mem_54[206]=8'h8b;
        mem_54[207]=8'h8a;
        mem_54[208]=8'h70;
        mem_54[209]=8'h3e;
        mem_54[210]=8'hb5;
        mem_54[211]=8'h66;
        mem_54[212]=8'h48;
        mem_54[213]=8'h3;
        mem_54[214]=8'hf6;
        mem_54[215]=8'he;
        mem_54[216]=8'h61;
        mem_54[217]=8'h35;
        mem_54[218]=8'h57;
        mem_54[219]=8'hb9;
        mem_54[220]=8'h86;
        mem_54[221]=8'hc1;
        mem_54[222]=8'h1d;
        mem_54[223]=8'h9e;
        mem_54[224]=8'he1;
        mem_54[225]=8'hf8;
        mem_54[226]=8'h98;
        mem_54[227]=8'h11;
        mem_54[228]=8'h69;
        mem_54[229]=8'hd9;
        mem_54[230]=8'h8e;
        mem_54[231]=8'h94;
        mem_54[232]=8'h9b;
        mem_54[233]=8'h1e;
        mem_54[234]=8'h87;
        mem_54[235]=8'he9;
        mem_54[236]=8'hce;
        mem_54[237]=8'h55;
        mem_54[238]=8'h28;
        mem_54[239]=8'hdf;
        mem_54[240]=8'h8c;
        mem_54[241]=8'ha1;
        mem_54[242]=8'h89;
        mem_54[243]=8'hd;
        mem_54[244]=8'hbf;
        mem_54[245]=8'he6;
        mem_54[246]=8'h42;
        mem_54[247]=8'h68;
        mem_54[248]=8'h41;
        mem_54[249]=8'h99;
        mem_54[250]=8'h2d;
        mem_54[251]=8'hf;
        mem_54[252]=8'hb0;
        mem_54[253]=8'h54;
        mem_54[254]=8'hbb;
        mem_54[255]=8'h16;
    end

    initial begin
        mem_55[0]=8'h63;
        mem_55[1]=8'h7c;
        mem_55[2]=8'h77;
        mem_55[3]=8'h7b;
        mem_55[4]=8'hf2;
        mem_55[5]=8'h6b;
        mem_55[6]=8'h6f;
        mem_55[7]=8'hc5;
        mem_55[8]=8'h30;
        mem_55[9]=8'h1;
        mem_55[10]=8'h67;
        mem_55[11]=8'h2b;
        mem_55[12]=8'hfe;
        mem_55[13]=8'hd7;
        mem_55[14]=8'hab;
        mem_55[15]=8'h76;
        mem_55[16]=8'hca;
        mem_55[17]=8'h82;
        mem_55[18]=8'hc9;
        mem_55[19]=8'h7d;
        mem_55[20]=8'hfa;
        mem_55[21]=8'h59;
        mem_55[22]=8'h47;
        mem_55[23]=8'hf0;
        mem_55[24]=8'had;
        mem_55[25]=8'hd4;
        mem_55[26]=8'ha2;
        mem_55[27]=8'haf;
        mem_55[28]=8'h9c;
        mem_55[29]=8'ha4;
        mem_55[30]=8'h72;
        mem_55[31]=8'hc0;
        mem_55[32]=8'hb7;
        mem_55[33]=8'hfd;
        mem_55[34]=8'h93;
        mem_55[35]=8'h26;
        mem_55[36]=8'h36;
        mem_55[37]=8'h3f;
        mem_55[38]=8'hf7;
        mem_55[39]=8'hcc;
        mem_55[40]=8'h34;
        mem_55[41]=8'ha5;
        mem_55[42]=8'he5;
        mem_55[43]=8'hf1;
        mem_55[44]=8'h71;
        mem_55[45]=8'hd8;
        mem_55[46]=8'h31;
        mem_55[47]=8'h15;
        mem_55[48]=8'h4;
        mem_55[49]=8'hc7;
        mem_55[50]=8'h23;
        mem_55[51]=8'hc3;
        mem_55[52]=8'h18;
        mem_55[53]=8'h96;
        mem_55[54]=8'h5;
        mem_55[55]=8'h9a;
        mem_55[56]=8'h7;
        mem_55[57]=8'h12;
        mem_55[58]=8'h80;
        mem_55[59]=8'he2;
        mem_55[60]=8'heb;
        mem_55[61]=8'h27;
        mem_55[62]=8'hb2;
        mem_55[63]=8'h75;
        mem_55[64]=8'h9;
        mem_55[65]=8'h83;
        mem_55[66]=8'h2c;
        mem_55[67]=8'h1a;
        mem_55[68]=8'h1b;
        mem_55[69]=8'h6e;
        mem_55[70]=8'h5a;
        mem_55[71]=8'ha0;
        mem_55[72]=8'h52;
        mem_55[73]=8'h3b;
        mem_55[74]=8'hd6;
        mem_55[75]=8'hb3;
        mem_55[76]=8'h29;
        mem_55[77]=8'he3;
        mem_55[78]=8'h2f;
        mem_55[79]=8'h84;
        mem_55[80]=8'h53;
        mem_55[81]=8'hd1;
        mem_55[82]=8'h0;
        mem_55[83]=8'hed;
        mem_55[84]=8'h20;
        mem_55[85]=8'hfc;
        mem_55[86]=8'hb1;
        mem_55[87]=8'h5b;
        mem_55[88]=8'h6a;
        mem_55[89]=8'hcb;
        mem_55[90]=8'hbe;
        mem_55[91]=8'h39;
        mem_55[92]=8'h4a;
        mem_55[93]=8'h4c;
        mem_55[94]=8'h58;
        mem_55[95]=8'hcf;
        mem_55[96]=8'hd0;
        mem_55[97]=8'hef;
        mem_55[98]=8'haa;
        mem_55[99]=8'hfb;
        mem_55[100]=8'h43;
        mem_55[101]=8'h4d;
        mem_55[102]=8'h33;
        mem_55[103]=8'h85;
        mem_55[104]=8'h45;
        mem_55[105]=8'hf9;
        mem_55[106]=8'h2;
        mem_55[107]=8'h7f;
        mem_55[108]=8'h50;
        mem_55[109]=8'h3c;
        mem_55[110]=8'h9f;
        mem_55[111]=8'ha8;
        mem_55[112]=8'h51;
        mem_55[113]=8'ha3;
        mem_55[114]=8'h40;
        mem_55[115]=8'h8f;
        mem_55[116]=8'h92;
        mem_55[117]=8'h9d;
        mem_55[118]=8'h38;
        mem_55[119]=8'hf5;
        mem_55[120]=8'hbc;
        mem_55[121]=8'hb6;
        mem_55[122]=8'hda;
        mem_55[123]=8'h21;
        mem_55[124]=8'h10;
        mem_55[125]=8'hff;
        mem_55[126]=8'hf3;
        mem_55[127]=8'hd2;
        mem_55[128]=8'hcd;
        mem_55[129]=8'hc;
        mem_55[130]=8'h13;
        mem_55[131]=8'hec;
        mem_55[132]=8'h5f;
        mem_55[133]=8'h97;
        mem_55[134]=8'h44;
        mem_55[135]=8'h17;
        mem_55[136]=8'hc4;
        mem_55[137]=8'ha7;
        mem_55[138]=8'h7e;
        mem_55[139]=8'h3d;
        mem_55[140]=8'h64;
        mem_55[141]=8'h5d;
        mem_55[142]=8'h19;
        mem_55[143]=8'h73;
        mem_55[144]=8'h60;
        mem_55[145]=8'h81;
        mem_55[146]=8'h4f;
        mem_55[147]=8'hdc;
        mem_55[148]=8'h22;
        mem_55[149]=8'h2a;
        mem_55[150]=8'h90;
        mem_55[151]=8'h88;
        mem_55[152]=8'h46;
        mem_55[153]=8'hee;
        mem_55[154]=8'hb8;
        mem_55[155]=8'h14;
        mem_55[156]=8'hde;
        mem_55[157]=8'h5e;
        mem_55[158]=8'hb;
        mem_55[159]=8'hdb;
        mem_55[160]=8'he0;
        mem_55[161]=8'h32;
        mem_55[162]=8'h3a;
        mem_55[163]=8'ha;
        mem_55[164]=8'h49;
        mem_55[165]=8'h6;
        mem_55[166]=8'h24;
        mem_55[167]=8'h5c;
        mem_55[168]=8'hc2;
        mem_55[169]=8'hd3;
        mem_55[170]=8'hac;
        mem_55[171]=8'h62;
        mem_55[172]=8'h91;
        mem_55[173]=8'h95;
        mem_55[174]=8'he4;
        mem_55[175]=8'h79;
        mem_55[176]=8'he7;
        mem_55[177]=8'hc8;
        mem_55[178]=8'h37;
        mem_55[179]=8'h6d;
        mem_55[180]=8'h8d;
        mem_55[181]=8'hd5;
        mem_55[182]=8'h4e;
        mem_55[183]=8'ha9;
        mem_55[184]=8'h6c;
        mem_55[185]=8'h56;
        mem_55[186]=8'hf4;
        mem_55[187]=8'hea;
        mem_55[188]=8'h65;
        mem_55[189]=8'h7a;
        mem_55[190]=8'hae;
        mem_55[191]=8'h8;
        mem_55[192]=8'hba;
        mem_55[193]=8'h78;
        mem_55[194]=8'h25;
        mem_55[195]=8'h2e;
        mem_55[196]=8'h1c;
        mem_55[197]=8'ha6;
        mem_55[198]=8'hb4;
        mem_55[199]=8'hc6;
        mem_55[200]=8'he8;
        mem_55[201]=8'hdd;
        mem_55[202]=8'h74;
        mem_55[203]=8'h1f;
        mem_55[204]=8'h4b;
        mem_55[205]=8'hbd;
        mem_55[206]=8'h8b;
        mem_55[207]=8'h8a;
        mem_55[208]=8'h70;
        mem_55[209]=8'h3e;
        mem_55[210]=8'hb5;
        mem_55[211]=8'h66;
        mem_55[212]=8'h48;
        mem_55[213]=8'h3;
        mem_55[214]=8'hf6;
        mem_55[215]=8'he;
        mem_55[216]=8'h61;
        mem_55[217]=8'h35;
        mem_55[218]=8'h57;
        mem_55[219]=8'hb9;
        mem_55[220]=8'h86;
        mem_55[221]=8'hc1;
        mem_55[222]=8'h1d;
        mem_55[223]=8'h9e;
        mem_55[224]=8'he1;
        mem_55[225]=8'hf8;
        mem_55[226]=8'h98;
        mem_55[227]=8'h11;
        mem_55[228]=8'h69;
        mem_55[229]=8'hd9;
        mem_55[230]=8'h8e;
        mem_55[231]=8'h94;
        mem_55[232]=8'h9b;
        mem_55[233]=8'h1e;
        mem_55[234]=8'h87;
        mem_55[235]=8'he9;
        mem_55[236]=8'hce;
        mem_55[237]=8'h55;
        mem_55[238]=8'h28;
        mem_55[239]=8'hdf;
        mem_55[240]=8'h8c;
        mem_55[241]=8'ha1;
        mem_55[242]=8'h89;
        mem_55[243]=8'hd;
        mem_55[244]=8'hbf;
        mem_55[245]=8'he6;
        mem_55[246]=8'h42;
        mem_55[247]=8'h68;
        mem_55[248]=8'h41;
        mem_55[249]=8'h99;
        mem_55[250]=8'h2d;
        mem_55[251]=8'hf;
        mem_55[252]=8'hb0;
        mem_55[253]=8'h54;
        mem_55[254]=8'hbb;
        mem_55[255]=8'h16;
    end

    initial begin
        mem_56[0]=8'h63;
        mem_56[1]=8'h7c;
        mem_56[2]=8'h77;
        mem_56[3]=8'h7b;
        mem_56[4]=8'hf2;
        mem_56[5]=8'h6b;
        mem_56[6]=8'h6f;
        mem_56[7]=8'hc5;
        mem_56[8]=8'h30;
        mem_56[9]=8'h1;
        mem_56[10]=8'h67;
        mem_56[11]=8'h2b;
        mem_56[12]=8'hfe;
        mem_56[13]=8'hd7;
        mem_56[14]=8'hab;
        mem_56[15]=8'h76;
        mem_56[16]=8'hca;
        mem_56[17]=8'h82;
        mem_56[18]=8'hc9;
        mem_56[19]=8'h7d;
        mem_56[20]=8'hfa;
        mem_56[21]=8'h59;
        mem_56[22]=8'h47;
        mem_56[23]=8'hf0;
        mem_56[24]=8'had;
        mem_56[25]=8'hd4;
        mem_56[26]=8'ha2;
        mem_56[27]=8'haf;
        mem_56[28]=8'h9c;
        mem_56[29]=8'ha4;
        mem_56[30]=8'h72;
        mem_56[31]=8'hc0;
        mem_56[32]=8'hb7;
        mem_56[33]=8'hfd;
        mem_56[34]=8'h93;
        mem_56[35]=8'h26;
        mem_56[36]=8'h36;
        mem_56[37]=8'h3f;
        mem_56[38]=8'hf7;
        mem_56[39]=8'hcc;
        mem_56[40]=8'h34;
        mem_56[41]=8'ha5;
        mem_56[42]=8'he5;
        mem_56[43]=8'hf1;
        mem_56[44]=8'h71;
        mem_56[45]=8'hd8;
        mem_56[46]=8'h31;
        mem_56[47]=8'h15;
        mem_56[48]=8'h4;
        mem_56[49]=8'hc7;
        mem_56[50]=8'h23;
        mem_56[51]=8'hc3;
        mem_56[52]=8'h18;
        mem_56[53]=8'h96;
        mem_56[54]=8'h5;
        mem_56[55]=8'h9a;
        mem_56[56]=8'h7;
        mem_56[57]=8'h12;
        mem_56[58]=8'h80;
        mem_56[59]=8'he2;
        mem_56[60]=8'heb;
        mem_56[61]=8'h27;
        mem_56[62]=8'hb2;
        mem_56[63]=8'h75;
        mem_56[64]=8'h9;
        mem_56[65]=8'h83;
        mem_56[66]=8'h2c;
        mem_56[67]=8'h1a;
        mem_56[68]=8'h1b;
        mem_56[69]=8'h6e;
        mem_56[70]=8'h5a;
        mem_56[71]=8'ha0;
        mem_56[72]=8'h52;
        mem_56[73]=8'h3b;
        mem_56[74]=8'hd6;
        mem_56[75]=8'hb3;
        mem_56[76]=8'h29;
        mem_56[77]=8'he3;
        mem_56[78]=8'h2f;
        mem_56[79]=8'h84;
        mem_56[80]=8'h53;
        mem_56[81]=8'hd1;
        mem_56[82]=8'h0;
        mem_56[83]=8'hed;
        mem_56[84]=8'h20;
        mem_56[85]=8'hfc;
        mem_56[86]=8'hb1;
        mem_56[87]=8'h5b;
        mem_56[88]=8'h6a;
        mem_56[89]=8'hcb;
        mem_56[90]=8'hbe;
        mem_56[91]=8'h39;
        mem_56[92]=8'h4a;
        mem_56[93]=8'h4c;
        mem_56[94]=8'h58;
        mem_56[95]=8'hcf;
        mem_56[96]=8'hd0;
        mem_56[97]=8'hef;
        mem_56[98]=8'haa;
        mem_56[99]=8'hfb;
        mem_56[100]=8'h43;
        mem_56[101]=8'h4d;
        mem_56[102]=8'h33;
        mem_56[103]=8'h85;
        mem_56[104]=8'h45;
        mem_56[105]=8'hf9;
        mem_56[106]=8'h2;
        mem_56[107]=8'h7f;
        mem_56[108]=8'h50;
        mem_56[109]=8'h3c;
        mem_56[110]=8'h9f;
        mem_56[111]=8'ha8;
        mem_56[112]=8'h51;
        mem_56[113]=8'ha3;
        mem_56[114]=8'h40;
        mem_56[115]=8'h8f;
        mem_56[116]=8'h92;
        mem_56[117]=8'h9d;
        mem_56[118]=8'h38;
        mem_56[119]=8'hf5;
        mem_56[120]=8'hbc;
        mem_56[121]=8'hb6;
        mem_56[122]=8'hda;
        mem_56[123]=8'h21;
        mem_56[124]=8'h10;
        mem_56[125]=8'hff;
        mem_56[126]=8'hf3;
        mem_56[127]=8'hd2;
        mem_56[128]=8'hcd;
        mem_56[129]=8'hc;
        mem_56[130]=8'h13;
        mem_56[131]=8'hec;
        mem_56[132]=8'h5f;
        mem_56[133]=8'h97;
        mem_56[134]=8'h44;
        mem_56[135]=8'h17;
        mem_56[136]=8'hc4;
        mem_56[137]=8'ha7;
        mem_56[138]=8'h7e;
        mem_56[139]=8'h3d;
        mem_56[140]=8'h64;
        mem_56[141]=8'h5d;
        mem_56[142]=8'h19;
        mem_56[143]=8'h73;
        mem_56[144]=8'h60;
        mem_56[145]=8'h81;
        mem_56[146]=8'h4f;
        mem_56[147]=8'hdc;
        mem_56[148]=8'h22;
        mem_56[149]=8'h2a;
        mem_56[150]=8'h90;
        mem_56[151]=8'h88;
        mem_56[152]=8'h46;
        mem_56[153]=8'hee;
        mem_56[154]=8'hb8;
        mem_56[155]=8'h14;
        mem_56[156]=8'hde;
        mem_56[157]=8'h5e;
        mem_56[158]=8'hb;
        mem_56[159]=8'hdb;
        mem_56[160]=8'he0;
        mem_56[161]=8'h32;
        mem_56[162]=8'h3a;
        mem_56[163]=8'ha;
        mem_56[164]=8'h49;
        mem_56[165]=8'h6;
        mem_56[166]=8'h24;
        mem_56[167]=8'h5c;
        mem_56[168]=8'hc2;
        mem_56[169]=8'hd3;
        mem_56[170]=8'hac;
        mem_56[171]=8'h62;
        mem_56[172]=8'h91;
        mem_56[173]=8'h95;
        mem_56[174]=8'he4;
        mem_56[175]=8'h79;
        mem_56[176]=8'he7;
        mem_56[177]=8'hc8;
        mem_56[178]=8'h37;
        mem_56[179]=8'h6d;
        mem_56[180]=8'h8d;
        mem_56[181]=8'hd5;
        mem_56[182]=8'h4e;
        mem_56[183]=8'ha9;
        mem_56[184]=8'h6c;
        mem_56[185]=8'h56;
        mem_56[186]=8'hf4;
        mem_56[187]=8'hea;
        mem_56[188]=8'h65;
        mem_56[189]=8'h7a;
        mem_56[190]=8'hae;
        mem_56[191]=8'h8;
        mem_56[192]=8'hba;
        mem_56[193]=8'h78;
        mem_56[194]=8'h25;
        mem_56[195]=8'h2e;
        mem_56[196]=8'h1c;
        mem_56[197]=8'ha6;
        mem_56[198]=8'hb4;
        mem_56[199]=8'hc6;
        mem_56[200]=8'he8;
        mem_56[201]=8'hdd;
        mem_56[202]=8'h74;
        mem_56[203]=8'h1f;
        mem_56[204]=8'h4b;
        mem_56[205]=8'hbd;
        mem_56[206]=8'h8b;
        mem_56[207]=8'h8a;
        mem_56[208]=8'h70;
        mem_56[209]=8'h3e;
        mem_56[210]=8'hb5;
        mem_56[211]=8'h66;
        mem_56[212]=8'h48;
        mem_56[213]=8'h3;
        mem_56[214]=8'hf6;
        mem_56[215]=8'he;
        mem_56[216]=8'h61;
        mem_56[217]=8'h35;
        mem_56[218]=8'h57;
        mem_56[219]=8'hb9;
        mem_56[220]=8'h86;
        mem_56[221]=8'hc1;
        mem_56[222]=8'h1d;
        mem_56[223]=8'h9e;
        mem_56[224]=8'he1;
        mem_56[225]=8'hf8;
        mem_56[226]=8'h98;
        mem_56[227]=8'h11;
        mem_56[228]=8'h69;
        mem_56[229]=8'hd9;
        mem_56[230]=8'h8e;
        mem_56[231]=8'h94;
        mem_56[232]=8'h9b;
        mem_56[233]=8'h1e;
        mem_56[234]=8'h87;
        mem_56[235]=8'he9;
        mem_56[236]=8'hce;
        mem_56[237]=8'h55;
        mem_56[238]=8'h28;
        mem_56[239]=8'hdf;
        mem_56[240]=8'h8c;
        mem_56[241]=8'ha1;
        mem_56[242]=8'h89;
        mem_56[243]=8'hd;
        mem_56[244]=8'hbf;
        mem_56[245]=8'he6;
        mem_56[246]=8'h42;
        mem_56[247]=8'h68;
        mem_56[248]=8'h41;
        mem_56[249]=8'h99;
        mem_56[250]=8'h2d;
        mem_56[251]=8'hf;
        mem_56[252]=8'hb0;
        mem_56[253]=8'h54;
        mem_56[254]=8'hbb;
        mem_56[255]=8'h16;
    end

    initial begin
        mem_57[0]=8'h63;
        mem_57[1]=8'h7c;
        mem_57[2]=8'h77;
        mem_57[3]=8'h7b;
        mem_57[4]=8'hf2;
        mem_57[5]=8'h6b;
        mem_57[6]=8'h6f;
        mem_57[7]=8'hc5;
        mem_57[8]=8'h30;
        mem_57[9]=8'h1;
        mem_57[10]=8'h67;
        mem_57[11]=8'h2b;
        mem_57[12]=8'hfe;
        mem_57[13]=8'hd7;
        mem_57[14]=8'hab;
        mem_57[15]=8'h76;
        mem_57[16]=8'hca;
        mem_57[17]=8'h82;
        mem_57[18]=8'hc9;
        mem_57[19]=8'h7d;
        mem_57[20]=8'hfa;
        mem_57[21]=8'h59;
        mem_57[22]=8'h47;
        mem_57[23]=8'hf0;
        mem_57[24]=8'had;
        mem_57[25]=8'hd4;
        mem_57[26]=8'ha2;
        mem_57[27]=8'haf;
        mem_57[28]=8'h9c;
        mem_57[29]=8'ha4;
        mem_57[30]=8'h72;
        mem_57[31]=8'hc0;
        mem_57[32]=8'hb7;
        mem_57[33]=8'hfd;
        mem_57[34]=8'h93;
        mem_57[35]=8'h26;
        mem_57[36]=8'h36;
        mem_57[37]=8'h3f;
        mem_57[38]=8'hf7;
        mem_57[39]=8'hcc;
        mem_57[40]=8'h34;
        mem_57[41]=8'ha5;
        mem_57[42]=8'he5;
        mem_57[43]=8'hf1;
        mem_57[44]=8'h71;
        mem_57[45]=8'hd8;
        mem_57[46]=8'h31;
        mem_57[47]=8'h15;
        mem_57[48]=8'h4;
        mem_57[49]=8'hc7;
        mem_57[50]=8'h23;
        mem_57[51]=8'hc3;
        mem_57[52]=8'h18;
        mem_57[53]=8'h96;
        mem_57[54]=8'h5;
        mem_57[55]=8'h9a;
        mem_57[56]=8'h7;
        mem_57[57]=8'h12;
        mem_57[58]=8'h80;
        mem_57[59]=8'he2;
        mem_57[60]=8'heb;
        mem_57[61]=8'h27;
        mem_57[62]=8'hb2;
        mem_57[63]=8'h75;
        mem_57[64]=8'h9;
        mem_57[65]=8'h83;
        mem_57[66]=8'h2c;
        mem_57[67]=8'h1a;
        mem_57[68]=8'h1b;
        mem_57[69]=8'h6e;
        mem_57[70]=8'h5a;
        mem_57[71]=8'ha0;
        mem_57[72]=8'h52;
        mem_57[73]=8'h3b;
        mem_57[74]=8'hd6;
        mem_57[75]=8'hb3;
        mem_57[76]=8'h29;
        mem_57[77]=8'he3;
        mem_57[78]=8'h2f;
        mem_57[79]=8'h84;
        mem_57[80]=8'h53;
        mem_57[81]=8'hd1;
        mem_57[82]=8'h0;
        mem_57[83]=8'hed;
        mem_57[84]=8'h20;
        mem_57[85]=8'hfc;
        mem_57[86]=8'hb1;
        mem_57[87]=8'h5b;
        mem_57[88]=8'h6a;
        mem_57[89]=8'hcb;
        mem_57[90]=8'hbe;
        mem_57[91]=8'h39;
        mem_57[92]=8'h4a;
        mem_57[93]=8'h4c;
        mem_57[94]=8'h58;
        mem_57[95]=8'hcf;
        mem_57[96]=8'hd0;
        mem_57[97]=8'hef;
        mem_57[98]=8'haa;
        mem_57[99]=8'hfb;
        mem_57[100]=8'h43;
        mem_57[101]=8'h4d;
        mem_57[102]=8'h33;
        mem_57[103]=8'h85;
        mem_57[104]=8'h45;
        mem_57[105]=8'hf9;
        mem_57[106]=8'h2;
        mem_57[107]=8'h7f;
        mem_57[108]=8'h50;
        mem_57[109]=8'h3c;
        mem_57[110]=8'h9f;
        mem_57[111]=8'ha8;
        mem_57[112]=8'h51;
        mem_57[113]=8'ha3;
        mem_57[114]=8'h40;
        mem_57[115]=8'h8f;
        mem_57[116]=8'h92;
        mem_57[117]=8'h9d;
        mem_57[118]=8'h38;
        mem_57[119]=8'hf5;
        mem_57[120]=8'hbc;
        mem_57[121]=8'hb6;
        mem_57[122]=8'hda;
        mem_57[123]=8'h21;
        mem_57[124]=8'h10;
        mem_57[125]=8'hff;
        mem_57[126]=8'hf3;
        mem_57[127]=8'hd2;
        mem_57[128]=8'hcd;
        mem_57[129]=8'hc;
        mem_57[130]=8'h13;
        mem_57[131]=8'hec;
        mem_57[132]=8'h5f;
        mem_57[133]=8'h97;
        mem_57[134]=8'h44;
        mem_57[135]=8'h17;
        mem_57[136]=8'hc4;
        mem_57[137]=8'ha7;
        mem_57[138]=8'h7e;
        mem_57[139]=8'h3d;
        mem_57[140]=8'h64;
        mem_57[141]=8'h5d;
        mem_57[142]=8'h19;
        mem_57[143]=8'h73;
        mem_57[144]=8'h60;
        mem_57[145]=8'h81;
        mem_57[146]=8'h4f;
        mem_57[147]=8'hdc;
        mem_57[148]=8'h22;
        mem_57[149]=8'h2a;
        mem_57[150]=8'h90;
        mem_57[151]=8'h88;
        mem_57[152]=8'h46;
        mem_57[153]=8'hee;
        mem_57[154]=8'hb8;
        mem_57[155]=8'h14;
        mem_57[156]=8'hde;
        mem_57[157]=8'h5e;
        mem_57[158]=8'hb;
        mem_57[159]=8'hdb;
        mem_57[160]=8'he0;
        mem_57[161]=8'h32;
        mem_57[162]=8'h3a;
        mem_57[163]=8'ha;
        mem_57[164]=8'h49;
        mem_57[165]=8'h6;
        mem_57[166]=8'h24;
        mem_57[167]=8'h5c;
        mem_57[168]=8'hc2;
        mem_57[169]=8'hd3;
        mem_57[170]=8'hac;
        mem_57[171]=8'h62;
        mem_57[172]=8'h91;
        mem_57[173]=8'h95;
        mem_57[174]=8'he4;
        mem_57[175]=8'h79;
        mem_57[176]=8'he7;
        mem_57[177]=8'hc8;
        mem_57[178]=8'h37;
        mem_57[179]=8'h6d;
        mem_57[180]=8'h8d;
        mem_57[181]=8'hd5;
        mem_57[182]=8'h4e;
        mem_57[183]=8'ha9;
        mem_57[184]=8'h6c;
        mem_57[185]=8'h56;
        mem_57[186]=8'hf4;
        mem_57[187]=8'hea;
        mem_57[188]=8'h65;
        mem_57[189]=8'h7a;
        mem_57[190]=8'hae;
        mem_57[191]=8'h8;
        mem_57[192]=8'hba;
        mem_57[193]=8'h78;
        mem_57[194]=8'h25;
        mem_57[195]=8'h2e;
        mem_57[196]=8'h1c;
        mem_57[197]=8'ha6;
        mem_57[198]=8'hb4;
        mem_57[199]=8'hc6;
        mem_57[200]=8'he8;
        mem_57[201]=8'hdd;
        mem_57[202]=8'h74;
        mem_57[203]=8'h1f;
        mem_57[204]=8'h4b;
        mem_57[205]=8'hbd;
        mem_57[206]=8'h8b;
        mem_57[207]=8'h8a;
        mem_57[208]=8'h70;
        mem_57[209]=8'h3e;
        mem_57[210]=8'hb5;
        mem_57[211]=8'h66;
        mem_57[212]=8'h48;
        mem_57[213]=8'h3;
        mem_57[214]=8'hf6;
        mem_57[215]=8'he;
        mem_57[216]=8'h61;
        mem_57[217]=8'h35;
        mem_57[218]=8'h57;
        mem_57[219]=8'hb9;
        mem_57[220]=8'h86;
        mem_57[221]=8'hc1;
        mem_57[222]=8'h1d;
        mem_57[223]=8'h9e;
        mem_57[224]=8'he1;
        mem_57[225]=8'hf8;
        mem_57[226]=8'h98;
        mem_57[227]=8'h11;
        mem_57[228]=8'h69;
        mem_57[229]=8'hd9;
        mem_57[230]=8'h8e;
        mem_57[231]=8'h94;
        mem_57[232]=8'h9b;
        mem_57[233]=8'h1e;
        mem_57[234]=8'h87;
        mem_57[235]=8'he9;
        mem_57[236]=8'hce;
        mem_57[237]=8'h55;
        mem_57[238]=8'h28;
        mem_57[239]=8'hdf;
        mem_57[240]=8'h8c;
        mem_57[241]=8'ha1;
        mem_57[242]=8'h89;
        mem_57[243]=8'hd;
        mem_57[244]=8'hbf;
        mem_57[245]=8'he6;
        mem_57[246]=8'h42;
        mem_57[247]=8'h68;
        mem_57[248]=8'h41;
        mem_57[249]=8'h99;
        mem_57[250]=8'h2d;
        mem_57[251]=8'hf;
        mem_57[252]=8'hb0;
        mem_57[253]=8'h54;
        mem_57[254]=8'hbb;
        mem_57[255]=8'h16;
    end

    // Combinational
    assign const_0_1 = 1;
    assign const_1_0 = 0;
    assign const_2_0 = 0;
    assign const_3_1 = 1;
    assign const_4_0 = 0;
    assign const_5_10 = 10;
    assign const_6_1 = 1;
    assign const_7_0 = 0;
    assign const_8_9 = 9;
    assign const_9_0 = 0;
    assign const_10_0 = 0;
    assign const_11_0 = 0;
    assign const_12_0 = 0;
    assign const_13_0 = 0;
    assign const_14_0 = 0;
    assign const_15_10 = 10;
    assign aes_ciphertext = tmp0;
    assign ready = tmp195;
    assign tmp13 = {tmp0[7], tmp0[6], tmp0[5], tmp0[4], tmp0[3], tmp0[2], tmp0[1], tmp0[0]};
    assign tmp14 = {tmp0[15], tmp0[14], tmp0[13], tmp0[12], tmp0[11], tmp0[10], tmp0[9], tmp0[8]};
    assign tmp15 = {tmp0[23], tmp0[22], tmp0[21], tmp0[20], tmp0[19], tmp0[18], tmp0[17], tmp0[16]};
    assign tmp16 = {tmp0[31], tmp0[30], tmp0[29], tmp0[28], tmp0[27], tmp0[26], tmp0[25], tmp0[24]};
    assign tmp17 = {tmp0[39], tmp0[38], tmp0[37], tmp0[36], tmp0[35], tmp0[34], tmp0[33], tmp0[32]};
    assign tmp18 = {tmp0[47], tmp0[46], tmp0[45], tmp0[44], tmp0[43], tmp0[42], tmp0[41], tmp0[40]};
    assign tmp19 = {tmp0[55], tmp0[54], tmp0[53], tmp0[52], tmp0[51], tmp0[50], tmp0[49], tmp0[48]};
    assign tmp20 = {tmp0[63], tmp0[62], tmp0[61], tmp0[60], tmp0[59], tmp0[58], tmp0[57], tmp0[56]};
    assign tmp21 = {tmp0[71], tmp0[70], tmp0[69], tmp0[68], tmp0[67], tmp0[66], tmp0[65], tmp0[64]};
    assign tmp22 = {tmp0[79], tmp0[78], tmp0[77], tmp0[76], tmp0[75], tmp0[74], tmp0[73], tmp0[72]};
    assign tmp23 = {tmp0[87], tmp0[86], tmp0[85], tmp0[84], tmp0[83], tmp0[82], tmp0[81], tmp0[80]};
    assign tmp24 = {tmp0[95], tmp0[94], tmp0[93], tmp0[92], tmp0[91], tmp0[90], tmp0[89], tmp0[88]};
    assign tmp25 = {tmp0[103], tmp0[102], tmp0[101], tmp0[100], tmp0[99], tmp0[98], tmp0[97], tmp0[96]};
    assign tmp26 = {tmp0[111], tmp0[110], tmp0[109], tmp0[108], tmp0[107], tmp0[106], tmp0[105], tmp0[104]};
    assign tmp27 = {tmp0[119], tmp0[118], tmp0[117], tmp0[116], tmp0[115], tmp0[114], tmp0[113], tmp0[112]};
    assign tmp28 = {tmp0[127], tmp0[126], tmp0[125], tmp0[124], tmp0[123], tmp0[122], tmp0[121], tmp0[120]};
    assign tmp45 = {tmp29, tmp30, tmp31, tmp32, tmp33, tmp34, tmp35, tmp36, tmp37, tmp38, tmp39, tmp40, tmp41, tmp42, tmp43, tmp44};
    assign tmp46 = {tmp45[7], tmp45[6], tmp45[5], tmp45[4], tmp45[3], tmp45[2], tmp45[1], tmp45[0]};
    assign tmp47 = {tmp45[15], tmp45[14], tmp45[13], tmp45[12], tmp45[11], tmp45[10], tmp45[9], tmp45[8]};
    assign tmp48 = {tmp45[23], tmp45[22], tmp45[21], tmp45[20], tmp45[19], tmp45[18], tmp45[17], tmp45[16]};
    assign tmp49 = {tmp45[31], tmp45[30], tmp45[29], tmp45[28], tmp45[27], tmp45[26], tmp45[25], tmp45[24]};
    assign tmp50 = {tmp45[39], tmp45[38], tmp45[37], tmp45[36], tmp45[35], tmp45[34], tmp45[33], tmp45[32]};
    assign tmp51 = {tmp45[47], tmp45[46], tmp45[45], tmp45[44], tmp45[43], tmp45[42], tmp45[41], tmp45[40]};
    assign tmp52 = {tmp45[55], tmp45[54], tmp45[53], tmp45[52], tmp45[51], tmp45[50], tmp45[49], tmp45[48]};
    assign tmp53 = {tmp45[63], tmp45[62], tmp45[61], tmp45[60], tmp45[59], tmp45[58], tmp45[57], tmp45[56]};
    assign tmp54 = {tmp45[71], tmp45[70], tmp45[69], tmp45[68], tmp45[67], tmp45[66], tmp45[65], tmp45[64]};
    assign tmp55 = {tmp45[79], tmp45[78], tmp45[77], tmp45[76], tmp45[75], tmp45[74], tmp45[73], tmp45[72]};
    assign tmp56 = {tmp45[87], tmp45[86], tmp45[85], tmp45[84], tmp45[83], tmp45[82], tmp45[81], tmp45[80]};
    assign tmp57 = {tmp45[95], tmp45[94], tmp45[93], tmp45[92], tmp45[91], tmp45[90], tmp45[89], tmp45[88]};
    assign tmp58 = {tmp45[103], tmp45[102], tmp45[101], tmp45[100], tmp45[99], tmp45[98], tmp45[97], tmp45[96]};
    assign tmp59 = {tmp45[111], tmp45[110], tmp45[109], tmp45[108], tmp45[107], tmp45[106], tmp45[105], tmp45[104]};
    assign tmp60 = {tmp45[119], tmp45[118], tmp45[117], tmp45[116], tmp45[115], tmp45[114], tmp45[113], tmp45[112]};
    assign tmp61 = {tmp45[127], tmp45[126], tmp45[125], tmp45[124], tmp45[123], tmp45[122], tmp45[121], tmp45[120]};
    assign tmp62 = {tmp61, tmp56, tmp51, tmp46, tmp57, tmp52, tmp47, tmp58, tmp53, tmp48, tmp59, tmp54, tmp49, tmp60, tmp55, tmp50};
    assign tmp63 = {tmp62[31], tmp62[30], tmp62[29], tmp62[28], tmp62[27], tmp62[26], tmp62[25], tmp62[24], tmp62[23], tmp62[22], tmp62[21], tmp62[20], tmp62[19], tmp62[18], tmp62[17], tmp62[16], tmp62[15], tmp62[14], tmp62[13], tmp62[12], tmp62[11], tmp62[10], tmp62[9], tmp62[8], tmp62[7], tmp62[6], tmp62[5], tmp62[4], tmp62[3], tmp62[2], tmp62[1], tmp62[0]};
    assign tmp64 = {tmp62[63], tmp62[62], tmp62[61], tmp62[60], tmp62[59], tmp62[58], tmp62[57], tmp62[56], tmp62[55], tmp62[54], tmp62[53], tmp62[52], tmp62[51], tmp62[50], tmp62[49], tmp62[48], tmp62[47], tmp62[46], tmp62[45], tmp62[44], tmp62[43], tmp62[42], tmp62[41], tmp62[40], tmp62[39], tmp62[38], tmp62[37], tmp62[36], tmp62[35], tmp62[34], tmp62[33], tmp62[32]};
    assign tmp65 = {tmp62[95], tmp62[94], tmp62[93], tmp62[92], tmp62[91], tmp62[90], tmp62[89], tmp62[88], tmp62[87], tmp62[86], tmp62[85], tmp62[84], tmp62[83], tmp62[82], tmp62[81], tmp62[80], tmp62[79], tmp62[78], tmp62[77], tmp62[76], tmp62[75], tmp62[74], tmp62[73], tmp62[72], tmp62[71], tmp62[70], tmp62[69], tmp62[68], tmp62[67], tmp62[66], tmp62[65], tmp62[64]};
    assign tmp66 = {tmp62[127], tmp62[126], tmp62[125], tmp62[124], tmp62[123], tmp62[122], tmp62[121], tmp62[120], tmp62[119], tmp62[118], tmp62[117], tmp62[116], tmp62[115], tmp62[114], tmp62[113], tmp62[112], tmp62[111], tmp62[110], tmp62[109], tmp62[108], tmp62[107], tmp62[106], tmp62[105], tmp62[104], tmp62[103], tmp62[102], tmp62[101], tmp62[100], tmp62[99], tmp62[98], tmp62[97], tmp62[96]};
    assign tmp67 = {tmp63[7], tmp63[6], tmp63[5], tmp63[4], tmp63[3], tmp63[2], tmp63[1], tmp63[0]};
    assign tmp68 = {tmp63[15], tmp63[14], tmp63[13], tmp63[12], tmp63[11], tmp63[10], tmp63[9], tmp63[8]};
    assign tmp69 = {tmp63[23], tmp63[22], tmp63[21], tmp63[20], tmp63[19], tmp63[18], tmp63[17], tmp63[16]};
    assign tmp70 = {tmp63[31], tmp63[30], tmp63[29], tmp63[28], tmp63[27], tmp63[26], tmp63[25], tmp63[24]};
    assign tmp72 = tmp71 ^ tmp68;
    assign tmp73 = tmp72 ^ tmp69;
    assign tmp75 = tmp73 ^ tmp74;
    assign tmp77 = tmp76 ^ tmp69;
    assign tmp78 = tmp77 ^ tmp70;
    assign tmp80 = tmp78 ^ tmp79;
    assign tmp82 = tmp81 ^ tmp70;
    assign tmp83 = tmp82 ^ tmp67;
    assign tmp85 = tmp83 ^ tmp84;
    assign tmp87 = tmp86 ^ tmp67;
    assign tmp88 = tmp87 ^ tmp68;
    assign tmp90 = tmp88 ^ tmp89;
    assign tmp91 = {tmp90, tmp85, tmp80, tmp75};
    assign tmp92 = {tmp64[7], tmp64[6], tmp64[5], tmp64[4], tmp64[3], tmp64[2], tmp64[1], tmp64[0]};
    assign tmp93 = {tmp64[15], tmp64[14], tmp64[13], tmp64[12], tmp64[11], tmp64[10], tmp64[9], tmp64[8]};
    assign tmp94 = {tmp64[23], tmp64[22], tmp64[21], tmp64[20], tmp64[19], tmp64[18], tmp64[17], tmp64[16]};
    assign tmp95 = {tmp64[31], tmp64[30], tmp64[29], tmp64[28], tmp64[27], tmp64[26], tmp64[25], tmp64[24]};
    assign tmp97 = tmp96 ^ tmp93;
    assign tmp98 = tmp97 ^ tmp94;
    assign tmp100 = tmp98 ^ tmp99;
    assign tmp102 = tmp101 ^ tmp94;
    assign tmp103 = tmp102 ^ tmp95;
    assign tmp105 = tmp103 ^ tmp104;
    assign tmp107 = tmp106 ^ tmp95;
    assign tmp108 = tmp107 ^ tmp92;
    assign tmp110 = tmp108 ^ tmp109;
    assign tmp112 = tmp111 ^ tmp92;
    assign tmp113 = tmp112 ^ tmp93;
    assign tmp115 = tmp113 ^ tmp114;
    assign tmp116 = {tmp115, tmp110, tmp105, tmp100};
    assign tmp117 = {tmp65[7], tmp65[6], tmp65[5], tmp65[4], tmp65[3], tmp65[2], tmp65[1], tmp65[0]};
    assign tmp118 = {tmp65[15], tmp65[14], tmp65[13], tmp65[12], tmp65[11], tmp65[10], tmp65[9], tmp65[8]};
    assign tmp119 = {tmp65[23], tmp65[22], tmp65[21], tmp65[20], tmp65[19], tmp65[18], tmp65[17], tmp65[16]};
    assign tmp120 = {tmp65[31], tmp65[30], tmp65[29], tmp65[28], tmp65[27], tmp65[26], tmp65[25], tmp65[24]};
    assign tmp122 = tmp121 ^ tmp118;
    assign tmp123 = tmp122 ^ tmp119;
    assign tmp125 = tmp123 ^ tmp124;
    assign tmp127 = tmp126 ^ tmp119;
    assign tmp128 = tmp127 ^ tmp120;
    assign tmp130 = tmp128 ^ tmp129;
    assign tmp132 = tmp131 ^ tmp120;
    assign tmp133 = tmp132 ^ tmp117;
    assign tmp135 = tmp133 ^ tmp134;
    assign tmp137 = tmp136 ^ tmp117;
    assign tmp138 = tmp137 ^ tmp118;
    assign tmp140 = tmp138 ^ tmp139;
    assign tmp141 = {tmp140, tmp135, tmp130, tmp125};
    assign tmp142 = {tmp66[7], tmp66[6], tmp66[5], tmp66[4], tmp66[3], tmp66[2], tmp66[1], tmp66[0]};
    assign tmp143 = {tmp66[15], tmp66[14], tmp66[13], tmp66[12], tmp66[11], tmp66[10], tmp66[9], tmp66[8]};
    assign tmp144 = {tmp66[23], tmp66[22], tmp66[21], tmp66[20], tmp66[19], tmp66[18], tmp66[17], tmp66[16]};
    assign tmp145 = {tmp66[31], tmp66[30], tmp66[29], tmp66[28], tmp66[27], tmp66[26], tmp66[25], tmp66[24]};
    assign tmp147 = tmp146 ^ tmp143;
    assign tmp148 = tmp147 ^ tmp144;
    assign tmp150 = tmp148 ^ tmp149;
    assign tmp152 = tmp151 ^ tmp144;
    assign tmp153 = tmp152 ^ tmp145;
    assign tmp155 = tmp153 ^ tmp154;
    assign tmp157 = tmp156 ^ tmp145;
    assign tmp158 = tmp157 ^ tmp142;
    assign tmp160 = tmp158 ^ tmp159;
    assign tmp162 = tmp161 ^ tmp142;
    assign tmp163 = tmp162 ^ tmp143;
    assign tmp165 = tmp163 ^ tmp164;
    assign tmp166 = {tmp165, tmp160, tmp155, tmp150};
    assign tmp167 = {tmp166, tmp141, tmp116, tmp91};
    assign tmp168 = {tmp1[31], tmp1[30], tmp1[29], tmp1[28], tmp1[27], tmp1[26], tmp1[25], tmp1[24], tmp1[23], tmp1[22], tmp1[21], tmp1[20], tmp1[19], tmp1[18], tmp1[17], tmp1[16], tmp1[15], tmp1[14], tmp1[13], tmp1[12], tmp1[11], tmp1[10], tmp1[9], tmp1[8], tmp1[7], tmp1[6], tmp1[5], tmp1[4], tmp1[3], tmp1[2], tmp1[1], tmp1[0]};
    assign tmp169 = {tmp1[63], tmp1[62], tmp1[61], tmp1[60], tmp1[59], tmp1[58], tmp1[57], tmp1[56], tmp1[55], tmp1[54], tmp1[53], tmp1[52], tmp1[51], tmp1[50], tmp1[49], tmp1[48], tmp1[47], tmp1[46], tmp1[45], tmp1[44], tmp1[43], tmp1[42], tmp1[41], tmp1[40], tmp1[39], tmp1[38], tmp1[37], tmp1[36], tmp1[35], tmp1[34], tmp1[33], tmp1[32]};
    assign tmp170 = {tmp1[95], tmp1[94], tmp1[93], tmp1[92], tmp1[91], tmp1[90], tmp1[89], tmp1[88], tmp1[87], tmp1[86], tmp1[85], tmp1[84], tmp1[83], tmp1[82], tmp1[81], tmp1[80], tmp1[79], tmp1[78], tmp1[77], tmp1[76], tmp1[75], tmp1[74], tmp1[73], tmp1[72], tmp1[71], tmp1[70], tmp1[69], tmp1[68], tmp1[67], tmp1[66], tmp1[65], tmp1[64]};
    assign tmp171 = {tmp1[127], tmp1[126], tmp1[125], tmp1[124], tmp1[123], tmp1[122], tmp1[121], tmp1[120], tmp1[119], tmp1[118], tmp1[117], tmp1[116], tmp1[115], tmp1[114], tmp1[113], tmp1[112], tmp1[111], tmp1[110], tmp1[109], tmp1[108], tmp1[107], tmp1[106], tmp1[105], tmp1[104], tmp1[103], tmp1[102], tmp1[101], tmp1[100], tmp1[99], tmp1[98], tmp1[97], tmp1[96]};
    assign tmp172 = {tmp168[7], tmp168[6], tmp168[5], tmp168[4], tmp168[3], tmp168[2], tmp168[1], tmp168[0]};
    assign tmp173 = {tmp168[15], tmp168[14], tmp168[13], tmp168[12], tmp168[11], tmp168[10], tmp168[9], tmp168[8]};
    assign tmp174 = {tmp168[23], tmp168[22], tmp168[21], tmp168[20], tmp168[19], tmp168[18], tmp168[17], tmp168[16]};
    assign tmp175 = {tmp168[31], tmp168[30], tmp168[29], tmp168[28], tmp168[27], tmp168[26], tmp168[25], tmp168[24]};
    assign tmp179 = {const_2_0, const_2_0, const_2_0, const_2_0};
    assign tmp180 = {tmp179, tmp202};
    assign tmp183 = tmp181 ^ tmp182;
    assign tmp187 = {tmp183, tmp184, tmp185, tmp186};
    assign tmp188 = tmp171 ^ tmp187;
    assign tmp189 = tmp188 ^ tmp170;
    assign tmp190 = tmp189 ^ tmp169;
    assign tmp191 = tmp190 ^ tmp168;
    assign tmp192 = {tmp188, tmp189, tmp190, tmp191};
    assign tmp193 = tmp243 ^ tmp233;
    assign tmp194 = reset == const_3_1;
    assign tmp195 = counter == const_5_10;
    assign tmp197 = tmp212 & tmp195;
    assign tmp200 = {const_7_0, const_7_0, const_7_0};
    assign tmp201 = {tmp200, const_6_1};
    assign tmp202 = counter + tmp201;
    assign tmp212 = ~tmp194;
    assign tmp215 = counter == const_8_9;
    assign tmp218 = tmp212 & tmp221;
    assign tmp219 = tmp218 & tmp215;
    assign tmp221 = ~tmp195;
    assign tmp223 = ~tmp215;
    assign tmp224 = tmp218 & tmp223;
    assign tmp226 = {tmp200, const_9_0};
    assign tmp227 = tmp194 ? const_4_0 : tmp226;
    assign tmp228 = tmp197 ? counter : tmp227;
    assign tmp229 = tmp218 ? tmp202 : tmp228;
    assign tmp230 = {const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0, const_12_0};
    assign tmp232 = tmp194 ? aes_key : tmp240;
    assign tmp233 = tmp218 ? tmp192 : tmp232;
    assign tmp234 = tmp194 ? tmp193 : tmp0;
    assign tmp235 = tmp197 ? tmp0 : tmp234;
    assign tmp236 = tmp218 ? tmp193 : tmp235;
    assign tmp237 = tmp194 ? aes_key : tmp1;
    assign tmp238 = tmp218 ? tmp192 : tmp237;
    assign tmp240 = {tmp230, const_13_0};
    assign tmp241 = tmp194 ? aes_plaintext : tmp240;
    assign tmp242 = tmp219 ? tmp62 : tmp241;
    assign tmp243 = tmp224 ? tmp167 : tmp242;

    // Registers
    always @(posedge clk)
    begin
        if (rst) begin
            counter <= 0;
            tmp0 <= 0;
            tmp1 <= 0;
        end
        else begin
            counter <= tmp229;
            tmp0 <= tmp236;
            tmp1 <= tmp238;
        end
    end

    // Memory mem_0: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp29 = mem_0[tmp28];

    // Memory mem_2: tmp6
    always @(posedge clk)
    begin
    end
    assign tmp182 = mem_2[tmp180];

    // Memory mem_3: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp71 = mem_3[tmp67];

    // Memory mem_4: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp74 = mem_4[tmp70];

    // Memory mem_9: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp30 = mem_9[tmp27];

    // Memory mem_10: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp31 = mem_10[tmp26];

    // Memory mem_11: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp32 = mem_11[tmp25];

    // Memory mem_12: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp33 = mem_12[tmp24];

    // Memory mem_13: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp34 = mem_13[tmp23];

    // Memory mem_14: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp35 = mem_14[tmp22];

    // Memory mem_15: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp36 = mem_15[tmp21];

    // Memory mem_16: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp37 = mem_16[tmp20];

    // Memory mem_17: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp38 = mem_17[tmp19];

    // Memory mem_18: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp39 = mem_18[tmp18];

    // Memory mem_19: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp40 = mem_19[tmp17];

    // Memory mem_20: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp41 = mem_20[tmp16];

    // Memory mem_21: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp42 = mem_21[tmp15];

    // Memory mem_22: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp43 = mem_22[tmp14];

    // Memory mem_23: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp44 = mem_23[tmp13];

    // Memory mem_24: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp76 = mem_24[tmp68];

    // Memory mem_25: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp79 = mem_25[tmp67];

    // Memory mem_26: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp81 = mem_26[tmp69];

    // Memory mem_27: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp84 = mem_27[tmp68];

    // Memory mem_28: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp86 = mem_28[tmp70];

    // Memory mem_29: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp89 = mem_29[tmp69];

    // Memory mem_30: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp96 = mem_30[tmp92];

    // Memory mem_31: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp99 = mem_31[tmp95];

    // Memory mem_32: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp101 = mem_32[tmp93];

    // Memory mem_33: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp104 = mem_33[tmp92];

    // Memory mem_34: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp106 = mem_34[tmp94];

    // Memory mem_35: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp109 = mem_35[tmp93];

    // Memory mem_36: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp111 = mem_36[tmp95];

    // Memory mem_37: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp114 = mem_37[tmp94];

    // Memory mem_38: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp121 = mem_38[tmp117];

    // Memory mem_39: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp124 = mem_39[tmp120];

    // Memory mem_40: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp126 = mem_40[tmp118];

    // Memory mem_41: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp129 = mem_41[tmp117];

    // Memory mem_42: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp131 = mem_42[tmp119];

    // Memory mem_43: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp134 = mem_43[tmp118];

    // Memory mem_44: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp136 = mem_44[tmp120];

    // Memory mem_45: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp139 = mem_45[tmp119];

    // Memory mem_46: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp146 = mem_46[tmp142];

    // Memory mem_47: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp149 = mem_47[tmp145];

    // Memory mem_48: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp151 = mem_48[tmp143];

    // Memory mem_49: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp154 = mem_49[tmp142];

    // Memory mem_50: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp156 = mem_50[tmp144];

    // Memory mem_51: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp159 = mem_51[tmp143];

    // Memory mem_52: tmp7
    always @(posedge clk)
    begin
    end
    assign tmp161 = mem_52[tmp145];

    // Memory mem_53: tmp8
    always @(posedge clk)
    begin
    end
    assign tmp164 = mem_53[tmp144];

    // Memory mem_54: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp181 = mem_54[tmp174];

    // Memory mem_55: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp184 = mem_55[tmp173];

    // Memory mem_56: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp185 = mem_56[tmp172];

    // Memory mem_57: tmp4
    always @(posedge clk)
    begin
    end
    assign tmp186 = mem_57[tmp175];

endmodule

