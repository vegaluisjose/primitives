module main(input clock, input reset, input [7:0] addr, output [7:0] data);

  wire [13:0] a;
  wire [15:0] d;

// RAMB18E2: 18K-bit Configurable Synchronous Block RAM
//           UltraScale
// Xilinx HDL Language Template, version 2020.2

(* LOC = "RAMB18_X0Y3", BEL = "RAMB18E2_U" *)
RAMB18E2 #(
   // CASCADE_ORDER_A, CASCADE_ORDER_B: "FIRST", "MIDDLE", "LAST", "NONE"
   .CASCADE_ORDER_A("NONE"),
   .CASCADE_ORDER_B("NONE"),
   // CLOCK_DOMAINS: "COMMON", "INDEPENDENT"
   .CLOCK_DOMAINS("INDEPENDENT"),
   // Collision check: "ALL", "GENERATE_X_ONLY", "NONE", "WARNING_ONLY"
   .SIM_COLLISION_CHECK("ALL"),
   // DOA_REG, DOB_REG: Optional output register (0, 1)
   .DOA_REG(0),
   .DOB_REG(0),
   // ENADDRENA/ENADDRENB: Address enable pin enable, "TRUE", "FALSE"
   .ENADDRENA("FALSE"),
   .ENADDRENB("FALSE"),
   // INITP_00 to INITP_07: Initial contents of parity memory array
   .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_00 to INIT_3F: Initial contents of data memory array
   .INIT_00(256'h00000000000000000000000000000000ffeeddccbbaa99887766554433221100),
   .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   // INIT_A, INIT_B: Initial values on output ports
   .INIT_A(18'h00000),
   .INIT_B(18'h00000),
   // Initialization File: RAM initialization file
   .INIT_FILE("NONE"),
   // Programmable Inversion Attributes: Specifies the use of the built-in programmable inversion
   .IS_CLKARDCLK_INVERTED(1'b0),
   .IS_CLKBWRCLK_INVERTED(1'b0),
   .IS_ENARDEN_INVERTED(1'b0),
   .IS_ENBWREN_INVERTED(1'b0),
   .IS_RSTRAMARSTRAM_INVERTED(1'b0),
   .IS_RSTRAMB_INVERTED(1'b0),
   .IS_RSTREGARSTREG_INVERTED(1'b0),
   .IS_RSTREGB_INVERTED(1'b0),
   // RDADDRCHANGE: Disable memory access when output value does not change ("TRUE", "FALSE")
   .RDADDRCHANGEA("FALSE"),
   .RDADDRCHANGEB("FALSE"),
   // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
   .READ_WIDTH_A(9),                                                                 // 0-9
   .READ_WIDTH_B(0),                                                                 // 0-9
   .WRITE_WIDTH_A(0),                                                                // 0-9
   .WRITE_WIDTH_B(0),                                                                // 0-9
   // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG", "REGCE")
   .RSTREG_PRIORITY_A("RSTREG"),
   .RSTREG_PRIORITY_B("RSTREG"),
   // SRVAL_A, SRVAL_B: Set/reset value for output
   .SRVAL_A(18'h00000),
   .SRVAL_B(18'h00000),
   // Sleep Async: Sleep function asynchronous or synchronous ("TRUE", "FALSE")
   .SLEEP_ASYNC("FALSE"),
   // WriteMode: "WRITE_FIRST", "NO_CHANGE", "READ_FIRST"
   .WRITE_MODE_A("NO_CHANGE"),
   .WRITE_MODE_B("NO_CHANGE")
)
RAMB18E2_inst (
   // Cascade Signals outputs: Multi-BRAM cascade signals
   .CASDOUTA(),               // 16-bit output: Port A cascade output data
   .CASDOUTB(),               // 16-bit output: Port B cascade output data
   .CASDOUTPA(),             // 2-bit output: Port A cascade output parity data
   .CASDOUTPB(),             // 2-bit output: Port B cascade output parity data
   // Port A Data outputs: Port A data
   .DOUTADOUT(d),             // 16-bit output: Port A data/LSB data
   .DOUTPADOUTP(),         // 2-bit output: Port A parity/LSB parity
   // Port B Data outputs: Port B data
   .DOUTBDOUT(),             // 16-bit output: Port B data/MSB data
   .DOUTPBDOUTP(),         // 2-bit output: Port B parity/MSB parity
   // Cascade Signals inputs: Multi-BRAM cascade signals
   .CASDIMUXA(1'b0),                  // 1-bit input: Port A input data (0=DINA, 1=CASDINA)
   .CASDIMUXB(1'b0),                  // 1-bit input: Port B input data (0=DINB, 1=CASDINB)
   .CASDINA(16'd0),                    // 16-bit input: Port A cascade input data
   .CASDINB(16'd0),                    // 16-bit input: Port B cascade input data
   .CASDINPA(2'd0),                   // 2-bit input: Port A cascade input parity data
   .CASDINPB(2'd0),                   // 2-bit input: Port B cascade input parity data
   .CASDOMUXA(1'b0),                  // 1-bit input: Port A unregistered data (0=BRAM data, 1=CASDINA)
   .CASDOMUXB(1'b0),                  // 1-bit input: Port B unregistered data (0=BRAM data, 1=CASDINB)
   .CASDOMUXEN_A(1'b0),               // 1-bit input: Port A unregistered output data enable
   .CASDOMUXEN_B(1'b0),               // 1-bit input: Port B unregistered output data enable
   .CASOREGIMUXA(1'b0),               // 1-bit input: Port A registered data (0=BRAM data, 1=CASDINA)
   .CASOREGIMUXB(1'b0),               // 1-bit input: Port B registered data (0=BRAM data, 1=CASDINB)
   .CASOREGIMUXEN_A(1'b0),            // 1-bit input: Port A registered output data enable
   .CASOREGIMUXEN_B(1'b0),            // 1-bit input: Port B registered output data enable
   // Port A Address/Control Signals inputs: Port A address and control signals
   .ADDRARDADDR(a),                   // 14-bit input: A/Read port address
   .ADDRENA(1'b0),                    // 1-bit input: Active-High A/Read port address enable
   .CLKARDCLK(clock),                  // 1-bit input: A/Read port clock
   .ENARDEN(1'b1),                    // 1-bit input: Port A enable/Read enable
   .REGCEAREGCE(1'b0),                // 1-bit input: Port A register enable/Register enable
   .RSTRAMARSTRAM(reset),              // 1-bit input: Port A set/reset
   .RSTREGARSTREG(reset),              // 1-bit input: Port A register set/reset
   .WEA(2'd0),                        // 2-bit input: Port A write enable
   // Port A Data inputs: Port A data
   .DINADIN(16'd0),                   // 16-bit input: Port A data/LSB data
   .DINPADINP(2'd0),                  // 2-bit input: Port A parity/LSB parity
   // Port B Address/Control Signals inputs: Port B address and control signals
   .ADDRBWRADDR(14'd0),         // 14-bit input: B/Write port address
   .ADDRENB(1'b0),                 // 1-bit input: Active-High B/Write port address enable
   .CLKBWRCLK(1'b0),             // 1-bit input: B/Write port clock
   .ENBWREN(1'b0),                 // 1-bit input: Port B enable/Write enable
   .REGCEB(1'b0),                   // 1-bit input: Port B register enable
   .RSTRAMB(1'b0),                 // 1-bit input: Port B set/reset
   .RSTREGB(1'b0),                 // 1-bit input: Port B register set/reset
   .SLEEP(1'b0),                     // 1-bit input: Sleep Mode
   .WEBWE(4'b0),                     // 4-bit input: Port B write enable/Write enable
   // Port B Data inputs: Port B data
   .DINBDIN(16'd0),                 // 16-bit input: Port B data/MSB data
   .DINPBDINP(2'd0)              // 2-bit input: Port B parity/MSB parity
);

   // End of RAMB18E2_inst instantiation

   assign a = {3'd0, addr, 3'd0};
   assign data = d[7:0];

endmodule
